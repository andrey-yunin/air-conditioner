��/  �}k�n��g,>�8����U$FU�R�H�� 9�Y�y�F�!�|o�-�ݨ��RAϪ�W�{6�!x�B��ux�v.5}�?UPݕ�O�#٤e��
��Z�޼�Cib"w�H�4_U,��W�^+79�������rc,�خ�bRޓ�+�|�O~g���!^�0d��o߹���ɯyw:=G�`�9�PyCE��8%X�7	]�*����pogU��(~X� ��Vrv����P�Uh:l���V�	�$���p�2��_1y�ȯ�u� 4�D�M��hݿDI� 6�pn�l�!`' ��-1�=<H_6�n�������@� ���Y�Q�`S-��O�Rd���pvTIuf���o?��q;���Ww�05�8)$P48�1z�j��=�j	���>Խ�ϒ�ƅm$oJY��Ғ<��o8?�8ƙ$6�@F�c�{�wah�$e�MwYL�2
��a��W���GN�R�#��O�pW�l�����Dꐿ&�~�i�w��Q�����&@q���}�s� L�]Z��q�TN��)��O���t`G�ev�bnl��N&�jQi��UX^2���e�%���&�2!"�}�2�zd
EJ3�0o>��u��b���6Ei�+^o�fr� �i��+��4����?�G���� ��M����IaeLMuI���4��ɪFG�sKRm۱������6������z����Y_ �����ޙ=b�*
[��L̛%x<ڵ����b�z`�.T�� ����Eݴ?��n��6���|�C�2p0�t�~�ątmOC�I'�.��D�ݧ�h�ȵ���<��@cW��'w�
����A���Vקr�y�3@�<؟=�Wo6u��BR��	o	���x�A����Ȏ;G9��cM��CW�e������2�Qr�.,�0l��xts�8�JP���#��!b�WC�A�MU@��P��nU�TW[�tVi�}���Dj/°�j��͓� �n-�ܹ�5d��[����Z_���y_W��T�b�@)�2�95��"��1:�[�R"�t�n,fw�9j�O�o�g0��,�!C�����E�TH���3�(V����W��LS���F�س��86�Z
a?0���uI����f�-��>�/a�zR6!Gp���zU�ա�{[D\��8?w�T�J��ӹ����
!'��r���;�S�&�szg@�I:�@^��\�l�J�0�y*�����-���qϣ�}2�A�yZ�]��k_YR�	2���̃�X����B��!v�J���ȐP�0�ğ���p��9��\?��
��TVe�O�k��1��V6��^8a���6V�TSiw:]���+���]�(i�&v�ܖ�³�)ش��&��0�:b�ý��1v���8I;,�z���;z����<�~��t�K��셐��lT�+��,�ҷ}�F���Mx{y��eT��`�a4�F��0�����+���=$.t����ԧ�U�g4�2�}�Z?�]E7D���ic�Wㄘ}��bN� _�O�K<X����߄� ��Чmw��X�`ߖ g���Y&y�&��]����o7N*b$ ������jW-1�{-�]߭�>Us;�c�3���7��ZfoQ��d08���%8��/s\�Z�\��Aq�R�5�M��z��I�SXh��IQ�|�e�f3� ����)ѥm��^��%CX=Km�I����be�M�E�m��+H��c�2��<�`���h�O��K�U�f�2j�����V�x0�����ɇ�i�0S� ,@��
�A�1���������&��w++�,�����]�7b������J� �[��<���r���>�Ka�0	n�V���8�KHuܽR&o��`2�(��FS�"�+_�:��ʿ����-�m �rG�S�V.�LP�í��;�F�@�T��WA�"�G*۟U�:��5pc�� �\�Kc���ǁ-L
Qn7w������4nO4�p�|&Y
�z*��0�'5�d_�B{�Aʡp�Y5��o36���2� �x���v+�"io��gv��V�J׷I.��n��x�h	s��U�S�*X7���T���rk�p�W-�;4�($��[�H���Hv}��[-T��>ra�2�Q��nWR�k񶢱�<�&��ho2"�3c�e��#��os���n�Ow�K}��|`�<nJԸ�Z�GCH�wzxF�4� ?�S�����r	N75�ʙ��'�OF��Q�_Ȳ����������[��G��u\�|}�U�׏�a��J����*>W�:�	��ߩN����t�Ub�����Dޖuj.�T�'W�f$J����Gl9��4��H��NU=�ܱ�=���`�V�	
6[@���I��8���d��g��.d&�(Wj	X$n7Ь���g\w\I��Dz��\58;���a4j�����O�0oo>�q\�5��]Z�L����L�Vuoa&����@7�����{��Nh�<���>��؛�=�J"�4;�q]g��c���ۏ��b5���	@l*�Dgc7�3�I��cȃ\��nIu�L$�!��O�8P�tۇ�''�����z��*�e}���Ⴝ�5�H�3"s�e�y��)߿G���
#h�Y�H����dq� (�zgY8��ۨ�3�@�I��A�����#Cd L�R�H�F�xa�gX���-��z�*�>�Ȩ�"��:L��:.�O.�Fj^���Ǒ�)�FF1f���f��^��	_n�M@4
+���$	�Ӛߴ/�ʌ�u�s�@����OMg�c��O�����U�2�ڋ�9��Б������;�����5U�)"d76?n%��$e=��"����c|M�8t�2f.j��W5\����V�DځL1��`O���J�H!��5r����!-p]u6K(�}��[����B�G�3�C�V���H<�G����vX�	�b�yxd��F
k�1�_'`L�*ɲ��$W��h'F�o�6��\��,��!�Ƭ9�Z2:����EƲ���+�oK��*Z��f.s�MI�����A��W������Θ�s2�t���m4�O;R(��LD�+$���+�nɭ���hT��k�y���+wn>x�k!Q���k)�F�J�`!	�d��w����L�`/�������l���9�����:�?�G��A�Ƭ�]��TW��,$� d�l/�κ��ì�;��
�"r �ip=��I���=YpF��}ӂ�.��--Ú#����0���#�6Y�J�ZN5��(]���nAn����Lh=�Ç 8Q�����CmW������S�;��>��<��p��D'_�31Uv����)�%U�Y��b��hJ"��;�Y3�ʰIm}���{�ֶG�Ƈ@���������E�zҊ���N�i�i�SpcΐT��/���D��h����&M���HQ�>�������O�q˂��(��RPh;�iC�_�a��s��H����NW`��k7��zm�ꑏ����4�T�n���k����!��zc��HNDUѶnz[XМrY(��j_}W] ,3; �p݋�>�5� �a�)n�n������6��(*�NM��#W�������GϚ ��R>B��Rc�	c�B.U;l�:�����[,�|��M��
f��rb<y��0d�%4[1h"#���i���(z׭�e���K(a��cRfo�-���|Z��s����X�,\ d|Ggi�*� :�4⛍F�!2�~�_*-�e��Y�y7��ū�K��_�[0X��Y?����C�Y���ܳq���2����!�F�w����-�(��&�I?`b(�����g$���H>���Hm��y�_�8N%�� ]�������_����IYe�B��eY·�;b_��?�IB�F"}ފoc��P0��g)Z�W��O��x}�{����Q4l�o:�����k�E�e�9�L��R�n1s��y��@�URD�F��󯬧�5A�h����4�'�4��(rR;��K:��.ѹ!�;�5[�nYZ�J�ŭ������j�M�ʔ4J�DE�"���sN>�+�m��d��5���К׏@�H���
�捷�ͽ��^'�����p{s"��%��?<�:�����k
q�c�Z�t!�?66߫d^���=m��m�5*R �8ڑM�s�L���|�|JEG��A�
nO��	��� ��پF�詰G[+���_��p��[���㐁6ç_�Ss�)�_���¤��kQXL��B^�BA���[ H�� ���H"y�3���ҟ�$~�~�G��v�Nۖ�	-·����:Y}���՘�>�#� �H��0:�9}JE����/����f����K� &��h%��Sh��ڐ�!a�o
��8�����:�Y�E����|�G-���i_��b���F*7��(T���ށd��l�x5�.���nS� ���8�_�,����G'��,
ufe3��7��o��,�y��d�n���Jd���% ��8�:�P�*I������.W�ӥ���}E�N� 7X���m�����%�,�~�J�ͫ$z����4 f��SzXTw��	Vh���ŴEo@����r��������.|��@�����P~�!  �_��������W��X59�Ѐ�N��e8lm!���۽��2�{H}��m#�+��y�1�NO��-���i�ZZdGC@@�.���H��
h��	��|w�V�c�LZ���k!�Q�k9}s�t{�c�v+f�����������HAjl�Yrz@KfѼ��������pW�B��wo0���{Q����63n��uB�c��7�a�	!+�,�F�,w�؞��80i�g���|��6$��� {��}�k�]1�(P�t,��}�֛��C1�;sou�"��ʪ'+cZ�o�P�bY*1�{;�����#�,��.�,!�P�����z!������9�wxIt蛲���?���N�G�&-����zP��g��`b_�����A� G�r.����!鳗�G:n0U;��}�jA����Z%��e� y�������,tnS��b�U����M��@��5`��>Y��7�H���h���I��(�qs��m�	Yה]��&����~�i��՚PۑMn�����":N�K 0�������lt:7��R�h�ů���Bw.�Ԥ,��(:/0��Ը[�!�~+���I.H�������z�V����i�2ԂȆr��6�<^:U'������ob8�J�����HB�ζ��*G+���g�[��2������(��⻓�sl�$��Y?��k�ө��`�v�n��"�c�"d+��K&k�U���O]'�-�碻�\��/*u�g:��`+ͱ;��k�a�y�P����}�}%�f��]��k�ҹ;��P�_���f.7��Z�9�He��p�Vd>�Wn�xYE0���u�H�(3����IC`Of=#�����L�P�\�k<㚄��6�#�:�Q/��Rq�:�NE�.��C/k�����"��p�E �_�I(R�U��EӾ~���LL>S��SŌ; o:x7Θ���3[{�����x�6�1�f-�P���uV��5�i�/2�M_����<��M�)�?C6X�Y���GbY���N���������V7�r��)��fF����FHjb@z���,�EOA4�5���a��f�g�T���N�<�M��$m@&��� S�<P� �u�ų[���r{�1r������)?�#���� ��x�J��Z�?X{+}�V0Q�N��i�&9E_&ߛ��]4�k���-�?:5uSQ]	FO�MR7�
��b�unydB~�C���+�_؍���a�wV�Pj���N�_$2K��uQ��I���--_�B>�|�/H.i�-q�E�+�W(��x�y�2ui�3S��ن�P�A���Mb������mQ*h�,���P��7!o��e������
al%�Y�� hP[��3Cn����˔[���Q��1G{�c�H`7�Y^��-8������3��~��$8��B����k�V�@q�5p�w۫[�*/�����]�nQ�OT����tv�B®n ���q��+����gf��HcL�U���<��D�j^����T����l@P�+��!T�ݦ�&o�4�@�eר�^���XΗ=���nUo><�E��F��(���G��
��.$]9q@*���O^Vd9vqvCDk-@��o�S����3���T�MY��"��f�Lm#e_$CF�~��B=�WJ���s���`:H�7�xF�/�&�p���M�:�;�MV����3ʃ��	q6&���d�w���8�ۜ$��\�G{1Q�n�$Q�i���2�5s���C"�oU��C������1�#'�2۴�/�!��(��� d	>�!j�oz�)�ae�
�H� ���}�*Yy�eUѠ�ԁ�~������߸�^�I���v�����i����}du���P�_Xk�Yϟ��+����tk�U�m������!$+�9�W؉�("2�D��ԇAʏ �ș�%�|�u/��� Ʌ�inzʳH�O��D ����]Pe:W�[ca�vv�l�u�<���] YHw��C�hfH�|Bzw{\L��R�m�F[Fv�1T�mPg|s�I�6$��>�E���P��
82R�U�w}����𜫒�iE 0|BF43͌H�}>�TS��Bp/xH��7o��4���gx�0c(�` � _����ٻ���OF�k���Vy=�QnZ|77�>�;�����JKS���BѣG-..�Фл��������}�����(�ݼk�^��3=R5t���䅜��]#��:+F�l_��x��⋷�蚚�c^/�,����al��Ng���7HP��V�>��4Wݢ���{���	,2Ĩ�<[���bt�<���+K����wLxGN�i:S�
\��q�OɈ&R�.���캳.�E����6���Z��"�gOu�ԯ��q����p[q�BHk�$��~� �0��Pᶃ8@k��;���^*���1�E^��� �E.{Mr�>U���ܖ��R7�h|��@�fK7����#Q8��?�_�s�����4�p�c�����-,�at@��	'���D+
�#{52[,��		t�`�dOX�����&o��1H��W9y}(�#GH�#B������<���ǫ�a�f#'��f��ȣ�(??[��7����Bˡ��_/п��wO�"2�i59k�ƺ�s[���ev֥��$jZ�����~�x��L^ TY[۱FL�o$�{i���ڀ�A�^�?4>�7, ���;�Z�M&n�u=���@���#�����C�:1�9�8P/���}���������&�5&����+*Eh��$�!�ADwh�C	J��-�6]���?z�jވc&w�P6hz�E��u���z�E߻P�1���fn������P�U��C����޳Z�'�E&}౦�"�)c����6����-�@E�|�a9�~TV�G�JM���=4{�hr���~���X�Vy~I�`Q��f3d��}+���y�Ͽ�7�X�)R��oq�R�^�z_�n��'�~�E�cu��Z�ܤ��d���5N�L��꤯�5ˏ<�n��J�+V�+�7�c�du/���z��̾#�L�����}�{�m�*��z7�A�������c�gج���5�ѝ��X� ���c ���a�(WW�
3��^�yK�R��rZw����bu�c'�tQ6��&}pt+��^;;\w���6�����f y���8$$�ktF?�q�9�����)a@TD���F\�]���<5��y�@Jha�ti�AI��/T-��G��$�y8rl�VD��;�S�Ո�O�~���N��ZsSFl��gj��Ӵb�W?\�6�bq
�(�3�������^DXC%o<�� )Y�qp��T�ĘD�1�$`�'^� _�
UK:�R�����:��vp�}gI�?`<4[��^��Nb���R�ќ����l��+$�qH�j��ꜱ���
4ʖ9SI��Ӝa�(�O����0������ƐL�R猔r�)Nhq��d̥�0wj��uI��f��Vx����nRm�x�OO��>:� ��쥞�ɹ�!����:���=u�[e��=b@��<P"yu��&_� �����ۋ?�9^mh08�2~��UχOoG�F�_��N���:�-[j��\?��(���o��)�䜙���G�����R�$�s�K	 e��pTe�"W^�2b&Fs�g�q��*��S�l�ERE�"Ec�ƪ������b�iR�y��#�@)��I�{�'�V?rt��x��Ơ��Z"X;r_��޶��A%K[�Z��ر��[;��U\Q������
1� 	n��'r%X��l	\o�st��(�Ч`�l誚��j[��·+�S��(R��^`wM͆dIaۃ-]B�׏��y-kBZ�ꖕɞ��X��x�Wsk���W"���.���l��@6�/���!3x�<��(LЊ�!�V��?4`��m��ֹ0�6����?�`��v]*�Ǚ��S�hf+�􃍄�/8�������(�7���M9��|����7&�G0�X^�j�]�����
��^�o��խ�<0}�`��)������6�+������NwA�J��\�~�5&��"	�[�	��5
� ����ص|�aLl�`s� ~��x%�#mã�X��=�,^sֿ�$�G;��c�VF�{� w��Y���ҍ�O��3�۾#������xE�*e�!�(��%�h���]E8�>#8�G7�ĵ롡	?c*M�L,���w@��htp��f2�C���C��e@db<T1�{&�%�nV�>d��5��IFc@�H��#��dJJzvы�*tM�iv��s��@Xa~Yc��dp���FF���.�K����Y'�����}�l�cI�Q0;��--w�� ���t��ۺ�~'�|�(j𷠤ǹ%���7"-��iG�:������K~�aLL��K)��Nw��~:��A����=;l�>� ��I�*`EQ���yI lUD �x�6����Ɖ�����uy�hs�c}Z��U`�v��ƅ�
�r)�ԯC��d�9a�G̵�=�����%�8�J�����2!�X�0�7L��lb1����>�@�O���$+�)���}7ٷX\�[*m�X���f�8݃-ڢʣ�