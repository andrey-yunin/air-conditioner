��/  �%��	����1�f���.m�{҅�8v~$�H���'Ⱉ��'�:7��բ����d{�nž@ɵoׯ�s~JE7�P����c������Q�R��.N�Ƶ�k����^_�#�ۃ�.Qz����ìF� Z�e�K����+qU�s�ލ�QC-���!^�0d��o߹���ɯyw:=G�`�9�PyCE��8%X�7	]�*����pogU��(~X� ��Vrv����P�Uh:l���V�	�$���p�2��_1y�ȯ�u� 4�D�M��hݿDI� 6�pn�l�!`' ��-1�=<H_6�n����X������y��I�����b�<W�Q�Ʌ�!$�;t�=��G�o�=�){�;Q���*%�8��P4�:�Ub�hQh�����_dzΎS@�׳�N4�$OO�������d^Q��u�ߪ[�C]�Y}N���*L���ql��~�F��<�E�!��=��=��~%�u���+�d�/bʾ(&fG/�����0j��k	��(����=�]4~�ŭ 侉����I2�_,,�g|3;�h���ԗ��HN�I�)��w�����ʮ�K.H��֌r��%��9��-��I��0�޾y�pTF�z]��l��1���0yoT�6Q�u�<����0 e�';�O���W뀬��f=��)���36�gaOnm��1#G�)L��T@ڀ|��][q��Q�	8��kp��S�ٿLyn��Χ�h�v���D}H+[@�Dɯ�7�i��+xli��r�.nǡ\i}`�ާ~N��.�#�t
[0��K�"'+��8(�bm��l�;�1���pr&sGR쨰������/�T��3ݙ~�y�i����)�Q�B&-���͉ �i�b�Qb�-���T���x@c�ȡ�r4�����5�a�#��B�;i���w�_e��"���H{�ơ3�l������\��w��K�H]������Dѧ�	��(ע��9��Kc;F���h�X/-�+���5XM3��=��3#����%��It���43�����1����,W��t��Y�.9¶P[���^��kȱ|�ߚ����7O�Ȁկ�����(�aR�7o�$���:�`�|���3e��w�	
��mI�B�۩����k�L�MG_�M���
ߵ	5��ݗa�F5�A�� 7��	(庺�X[~�����0�R��e�*��o�s9�B�EN�kq_ι����piZ_�y���
:�8�b���W�w8�Յ4G~(O�xzm��]v*��E���T�@O����U2�f�%ʩj"+�(Z���㜟C���;!���w�h�b�'v�q]}R>�͞Z���*�m4��P|���) �� �dOm)tX1���� R��Ġ=��H<X�"��t�w��=����m�V>�d������6�+��L�����ՈBk��|�F����f�'�+$!�����ޜyT*=	�J�{�/Ij�J)����YdG� è�N�~����썵׳~T:d�2Td5������n�,���E����E�|�/�nu"o�L�ɨ{�`;���#s�z�>*�U�1<�}}@�?6�m��A�&dS(�C#gv�\���k!,��)/�2m[�X�ք�,�ЯҮ��Ԓ�P
(a��z�(��Ga�Ɵr
b��si2�_�Mc�"~o��o֡l��)R4�'��AI�X�#�h6
���^�a��2ŀր���>�۝�cr�_bd^��Wr\�JX�h����:��@��3�y|�0h�^Gt��c��,E4j���paWY ��huJ
�'u�Im춋�;�vJƼ6�Hx⿎'׍���ܾ7f��Ȫ����m�V�b:rC�#�1��rت#6�,��c��A�޿w?D�ҷj�UǓ:+~�M� +�~*��K麆vSU�w��)Gw�Մ�n���7�EF��X^��e cN��-�D��k#U�
e�g~E��BV!�&�k�.���v�Ї �:�}B�_ ��ӉeKO[��α6$����[p��HM&x9j�M�
���c��,|�A�>2��9n��#��ǲA<U���NA�&&�D!��Bfa#"k�8�e�<)M����_�q+�/�612�+4( ���l�S8Z+r=�%>0J�T+�4����U�tٹT#[��J�ѯ��s��t����R�Bap���!R}Ƴ�qc&c���升r�fb+�!�E+��n�^��%RA��*�=���J�HIoQE�6���DO�bk-P������)�h{#�� ����o�Ll�+
sYf'��z9y!����Xʰt���<V�w������[���m���';l)~~����ijn�U��\0���O��e�o�n�� ( n����^D �ĂΖ�ۭ*�c�k�c���B������K�%`����J��|_��X��!�}xCH%�6�J�v]��p-���Q/;����	I�ɶz�4�e� _-��1���@��%���E�S�+�,�59]�q�?�%mUAǫ@@��д��=�Q)�x��&���-�#��>�bY�ҹ��
xj�T����'�_�4�W�+�:@�R�\�rn�Yz���Q��ռ�-q�R�Uő���4�Z������ �$e��e ��g=;�Lh�l�`:���KwJ3�α��s�lgH1-���+e�wm�>����4�c��)��V:�X�]ۗ0����-��UJy�����Gd�}+��l�;fsp �Mj?�����>yqW[�ss��xi��w���OB��˞1�����)�(�;[���Z/ ���P�S)\֢ON�aG�rS�����~���b�3΢YW��B{nd��AQN�O�Z�! �̄�)�9��<�Wj���z���r|���p���5��l��V��^�Q�!�NR���O�I��3�� �
���˘߽D ��ɿ?��ȯ�#HF��n���9z��!��Ĵ'���z\4��	��E�T���CDl��4MרƦ������n,CNW_��&
��g�V�yK�|�L}�V�Ш��cѿ��sD /h�r$0���4��ni"�dD��!��?���ȃɣ1.Y���5\�ֳ�ҟub���ϡC��C=~v�ߌ�x��,��+���z�q�1�J�E��w�H7A�&�"݉��ss�G{��i� >��jY&s��}ϧ���U����J�w��;n��"��O�iFݘ5B����X���@̰�(+P/�O�g*�z�_�[�2���ߢu���a��K�Ϫ��lv�a�����D��2�>Pj���:d�?c��zx������z^�����$'m7Ki�g|�����eB�ڜDG���HE[�AGB�>�L��kN����%Z�"�u�j\WF�'K7GvE�M.���ܱ��ٍ�kXdnU�t�n���q�b&C��g����S�K��r6q��r%"��#��~w>�(�����½�.��Ț��靈��Jw��3[&���	(�<aL��Nf�5��"�B�Լ�j��v���v����B�����;�~��h������̟�d��ں�r|�W�k���_���O�55l�b�/d��Fa���S|�e]�t�ē��g@�������g�압;��U�	󪜴�u}�n��)�6H�tǼ	�:c��ܝ�������]/M5瓓���`��(��i�|ї�FZ��x�5��}����Q)&p&abl3,�|����KJ�����������碘���ܓ�YeJ�;
��bݐ���4��~&zmY;�ȸ�+��K'�0Tn�$��Y&֪Xi4҇7�՜!\�BnL�C�(J ��������B :��!d� �{NB9������V�x ���T�̀�+�ӳ��d���bm{Lpþ!A~��� _�VO����e�2��k�y`�df�q &&����B.4�����6Q�E{���&-�3�⺍�fP�
�d�jA�����)���|�`�\��������j��(���¹$ Շw���=l�xL=v�����������#�K��?�D�?$���'t6X�"����e/�T��qv�=l�H�zC\`p&��R����1#����~܍�Iw�!o����!B�ڛ���6��b��_��{���fU����ݏ'���f�����s<.�Ň?���7����Qm�섊���w����l��A��j�7�9���H����ĳB��FJhy�&��Ƚ W�⃔�,�_�u�0L2�4�Q@�.��k����ub�"��
v�QV4ϴȲŲK�{�Tx2ՖNX�H�u�m�񵹛�p`~�e��]��=%��=��gi�U��&����f�3�����#�\H�C'�I��>Dh}B=��|�:�C#4 s�Ո���&㥩j�Ɗ���g�IH�1k��m�y�&pR9�(���K��8$$�c�P���,$@rm���➩���(bcV��n �C�|�o1���7�XMD�y1+���EWq�l��L�8�&}��b�>Ů5���y����vM	sc~j�F�`u��<8��[�i�LH5)�zP��Bnyx�r��/ )����-D?'K��_t���C
��3�2����7���Z��=��`*�4w����7�� ��VT�)�1rԬ��`��	�e����D�����LWgK�b��8�dgd��n1�Z0�,�6s��� ����b�$Śk�D>�q9���o�h���C/��7�:��� ��M��H��i�5��,GGQ$���t~��[?p�Zf�/FgW���cz�dۂǽ��Z�/qe|j���_���y���_�X���PK�<�ݙ�&�I�������k���v�?�O]Ř��भ��qN )xq��W�����!�R�ݧD�WY!m�ܧ�C��i�~�u���-�үξ)7�d�f�$i(tQd�|�\�r(�;�Uaye�p�&�.:,=�y+����t���1��1̓!9� ��/{Odg��9R\�q7� 8v����M�tk���)�d���E�4M���O�N��[�{u�tAS��t��� ��a�@_a8u�'z]yZ~�_�
�_,�.$L�ٻ�觙	�@�/m��p��uD��d��h=�/]������E�_Q]M��'N�r�b1(�G���-[Pe;Z+�+���-v�B_��������b�OOTM'_��~\2���Qo���}�\3��K���)!d�8�I��V��B�΍s6�p��U�2Y�����>�,2]R��~��,ܗ��e���&`f�^Yz!��� �G�lJ�>?�H2��5�Olp����w�[<3��G�I[�fȼ�>H@�F�L�+n��9��^�����@�ʔ �Β5�m�o�9lYHݢ<w�ps�D�,�6&VT�рo�n)�xĎ_F��_,��f|��!���Q���+	]�*��l����;�3�x��ҵ���ƙ��m��@(�ۻ��C]���_�U���A:usf�M���"S��f������ �1�����z�[�?Чjg��$������d��͝�'ψd�ݯE��g�DfR�m.�������#ԅ���4�WC-��.�j>�6xf�]+�u�tUU��(+�~�o^p
~�?�N����G�.����('�F6a�g?�H?��+�{cAt�rv�ɪ�ו@�p@v�Nm��7on6�����eyG������vw4_!��)y�� �$*��&=� *zfy�K��}�:\ֽi��w1ӭ�kk����tD�57Q�7��G��;��שމT-��Nh.^5fcC�e��H�p�����]�b&RC"���˃��9��L7ܘ;V��+'�n�?�[.��:�k+A�np�g�I�O��)=\��u��d5a�"y�&n7�gQi5|]D�z�4�y<�Z�Z�j��ى!�S��q��@lT�"�|�O��Q��P}}A�R#�.~��8�ꄺ�p�z�6ˤ�(���"��N��Z�w�a[Y��it��)��	�a{GF�h�@���btPvD%�e&��B������	�(Jڇ�{��Y�~Y6�Ag��N��[��{(y��Y��iw�h4�9���z#�K��K�@�վ4�����"�,�.�(�OF�No_��)�����������y�D�	��٣�g\:�w�
�SM2ŤqɪR!���Wol����a��Xl�����`l�gBa���X���\�\�wС����	%�R��c���|��D�A/�t��&��iܚ�~1�5�.�_,:�׈x����4i��Í7�1$S����4����̇�x��q���]�zѿ���LⵀH���kA^�$����w#�4�N~V>y���fok�}6e���g��;=c�yЇ��;-���t�g"��l�6������!\ ��.�OSqL�|���1�D@�{�@A򯱍ϥ�$Cr�R�C�L����,��-ByBFl���U�]��_�8*��ZB���?���"%�V��~�����l��1�CJ�J;���c���|ö����Tq\w�g�c��~������ى�IVA��g��<l=ZlZm2�I��w2���(8mfJ�a�g��ۯ  ?����C\��اϾM_��r,K"������'�y)b�Cs��]�C�.����PJ?�6M�$���5�3;±���������(u���!uqR��&�7�I4{@8��/A�D��y�-���$��V�B�I|ʾI�En�ub�n�$�*fw��\6��hU`gjL�x
k�Q���Ee+�Wh�$D=X��
y|pa���������嵁{���0�X,���.��*e��p���w���1�s$�{ۊh <�QZyO�=�t����_�LmHI�8�k_����3�1��Z@�p@?�n ��p6�'8�ÅgGӧ�y�c��ʄ��� {%r<����z6�����E�zM�Y\0j�>:�lӢS��Ӵy���@+�s6U��}����;����p`����;�<D/�Cr_ �xu (��V��W� ��NG��97:�ޔ���W���`�Mk�����J�W�El;�OA���D�L�?ф�LU$8�ґ����h�i��!�`�3}I�U"T뼑�����vB��*�z�J\k/l�D�X)b�F���)@%�����k��Kt�z��پ���7�,On�`��.ivM�HXgڗ�{i,��;o��y���J򣠅����ݴ^��{�ZV�!����ٯ<7/���{B%E���46�&zNZ��\��K�`W��;��c���E��S%�:Bm��=���]"�h�e�٘6����͖�����fmR�ƽ�o�V�j���&��lǪ@�!_���?BݲN!C��P`�	c���'�E׊ϓL��x��	�j_�_�$����Pߕ��mӤN��]�S{y^/>��	R�6�s�.ו�.7+�d{M8v�~1E>��e�B�����:�\��f�ka{�I�:���Q�2Ϲ�lԚ=�^6��lH�;Q��/P�`�8����[=^�PXls�(mYJ�C�;����a���[�	m��1�wd��L2�;M�-����@��l�i.?�VtGg�� �\C)�(m��K�ӢL��ZA|L�)�z�k�Ǳ�Ϫ�x3�J�8�Rc^û�6��)��	v���y��WRh,��.P5�9��c��s�=�f#u������P� ���uQj�����4)@TH�vV���\:�U�k�E~0W�������$ T]�>E������=�k��cd颰���,�����Y�����s^S�]�]w�*!�w���'�c�b��;sV�26ƒ�\	ց{S��,˃}�QT�;� j7s��-�o9�/�yg��`��1+r>�]1T��$����_�����E�t�Q1X	6�*!�A�g��`��7�pj��A�~CUXx�-����jȭ�.�������Ĺ�l��^4|�6R �h���p�LI�vU�_�Vޫ���Z}r�5��t��.�A�u�}ҹ"�yP�ÂE`�kj#�jj��j8�f׮�O���&�D�[��n�U
/B�P�V���p怊��-<?!%�B;�ڛ��B�u�]�B�F�3�o2r>>	��L�<B�{#O��1���$�At��T��\�ݝ����8����iA��BU�ʫ��S�&]U�3�ؖ��eW������yer���j����9�~f!�W5��n��T�n}r�߭ެ5$�I`fm̰���T��afGkʴ��8
���H�6��v�I=}61���:ºv�U,�6/�;bxw)u��W��G{`���I{M�^�a�-� ]��'#�Bu�!}�	~�-�Ȍn�1�i6��غ" �t���&�MX/�&:�ߕ���O�3v��|tj�ն��ЂH� X�/����>�U���t�tB�蚔����ݚ^5��x���,��ǚ���<\�� �Hm;����HoT/�AX�԰Q�W�Jό[R���n�ۍ#Uѹ�0� j.���>>�د h>(��Q\�
X�>�)��i�*n-ɷ��;��̵��I��D�E0Eʵ�5�������6�4:�sF�����)��x|��j��'�;����<�\�4����篘|�Ǳ�/4�+73v�\;�����P#����j�n�qG+������د�@�-�pw���(��/������ �B�c\v�Mh�f�[�?�5�i��/�"�tE.9a!�2k�y��/<>�� �RM��X�P�K={3��r�(�����_��B��J��$�"!4 
e-��c�*`�h3�uԚߑ��m��Gg�xv� �Њ�pg�SJ��yL�:��w�r�^GԞ�ԅ�#'ac˲��P�'s>F� P��o;��ˤ]�ɝsm���í��F)F��.}L�[A�Ҭ����w��!�����#}'��"��C52���H?9�m"@H���d�M:5�O�Rs���F&/�^n��ܭN�-0a����Ϻ-i*3��s�B!�jw�A�٥F���ǁ� Gv�:��&%�:멕��=���@]s�n9q:]���H��㸵>U ��0�����@�7���.�DA�O��G�A���.�|�z�4�~�F�물*� �X_�#d�_���A��O�#�9�Òv�URQ
�œ�
z鹘�̅(�e� ������ﵞ�ȼ�y��M��ѭ�f�<�3��,3<M@�J)�'����������;�E�>ޅEo����Ъ���V�O\�"xH���ȟ�2��U$-`H��)�Ͳ���]g�~�(r�KuY��MD�8׵T�T��dY�d_���C.�W���tb�HX<|e�M�or-Da�AK%:�w�Ԕy.�� �Y|tl��%�78k�� Z?Dc� �V��L)��J�|����6���@��>ͻ��-|�#
�����w��!���J���'����ٖS���1ӛ�����]MđH��H��:T�ܥ���#�ٻ����'uӇ��"�:�����s��{�MҪp>-MX��LvKE0fk��>x�4�\]~�U��8�ƧM��="�ŗ��	�c^u��9��O_U.�"N���ꛤ ;.�*K��zcv:a�b�є�%��VrP��T�vr�\�_g$�h��m˃������K�^ �BWI���K����b�ӳ�G��Xg�R4B
��eM�|d�'�y~���u��f��7�#��-�m�W3����pNn�f��]Y?�T�~���~����(Z���tU,tA�P]��-��:��з�SN�8rU�V���l��u�����͠�]3��t��Afu��:s�éq�k�<b�^��*vQ�hdI�t�V�����_^N�Jϻ;��M*9�*��c{�6�XqE��g6�Í���1��4X��Ǉ+��V|��1�w�h	��u�e�x�Ao{ޤ\�ߠ�_��G��&6i�!ڞ"���Zd.U,y��O
�#Th�Ū�%1�!��kB�&��8Y��,�	.��	R�np�A�!�K�G��:>J�f�s��܍�z���"p��Zm�P�0�d}+��F���&�?s�\��(���l^�s�sؔN-1^��Kp��XT(r�,3�j��ϯ�|��Vٸ�5�b&�PT6�Z��֡�t����i�����i0����5�%<��IԱ�2��#q̝8L��K V��byJ��t���QPS���4�6��>`|�$�n�S�\��U�S�`#������Q��*��%8s��X�p̉��MѢܢ������V�C���+~(�az�9F��?#����)�hC��Z�P��G�:�o��v�2%�~�����w���T�E�~��	�|>�zx��C?$��J뷧�͌�5\�3N�J���~���S]�Dw���!h�}�����+�ã+l�1�Q��w�Q���3�d���"aW�.�f�.��ww��5���>.s�)��嬚Cl��:ż�ٻ�[�*Q
y�¤���~/-$��X�� ���-6c�\Qj^G��T1��ٜY%��XqB�P�@<�ǖ����m��ȔD�5`�}��Z������Q,n����]�q^��rJ�]:�X슢�>c,z~#�������^`.�U�f�x�y��o����ǿl.7��X����Uո��ާ���>�H�Iٍ���}����P��w�Xz�6�-�A�o�
;�[Jv�l�F� Ds]=�Ͽ�n��^&�l$H�m��=꒮��c��������_a CU�3�s{n�J�4f}d��p7#.mn?� �iEC�f>{p�9ӄC�bʅF�lt;~Z~�+.ͬP�k/�2��wm�H��+��cÖ���* �I��ݯ��Y��^�{��]O3b���R|�]��
���m���k�I�iQ�6"��<����=;y�(� `)�):
�<
�����m�'d+�[yr�?����1� [ _Ԗ�`�D�
���r�8!��f\tc�,�E��r��:z�c�����|��	����4RR��~L x���mB쬞M}V���Ӱ�(��׃��7%rv;^_k��<d�̼���ܒ�@d!��� �����>t������7#Y�X�O]�}�oq"!<�y3$�1(�Y��޴ ��K��	�3]�Q{�c~;qj̓XE�~�1\o�������O:���_�H��FE����(�iG��d�k���"�И��/��v?��9���7�V�7�Mp�xŇ�jԺX�G�WL?��v��|��7��b�й	�'�.5n����bP�<�d00�;����7��J��K)f��T�p�\cVl#$�o��xt��,��c��4Q�-=}�x��Ê����1��`D�ٟ}������a���<ސ¶���u���"��~�P�xWS?��U_Q�e�<�� �e9�J�[=wCm\��9q�Z:{���z�s"����(;[��/�5�3��KVu��	J���u��[�8�������M�>kE3�z,�tK]��0�JLZ�裡[Mq�t�bB�8Y����4�A����;�+�W�/����pi���6���=R�ȸy�8g�_Zɱ��!�d�2��:���(�R�d�]e��{��J�b|�ڱ 4��&Ӄ��l�|�nPX�M�^�L��v?��c����u�"����yA��)���n����
N�UA����`���G~�Ih7�J�(���xN�<�Z�,���*:5gQ�&P�#φ�p��U0�,8�߀�ip�B���9ýI��DUeF��Cd>7w���L�~�L	}\f�)Vm�����N��I2�y��|J��~dP�=�Ms�����-G^>�͏�*`d.�h�7�j�_O�?�Xq��K]9�m]�ɓi�$��/ז�WFf��DWЉ�z��K��Z��hr�C�����m�ۧ��v��8�}����f�� ��2�'O��Ș��4��u\E9}x����,C$~����dq9-�,@���@�-]�ߎL�vM���K!�SС�`
F󿰢�%e���Z��~�t���]�����m!4vJ�������F��CC�Ȳ[��i�1HEb$6R��d��1=����/���6�����Э� e��R���M�Z�t|5Vuc�>��	����7�������3�qEl2�X���Y`5��k��e��]$�hRQ��S�S�t�;ĳڶ��6����Mt��o	ة�p�ѳ���v�W���`��,o�0^�1��&p������Qe2���q����f�An%tҿ���A�p������6��9�\%b���݇�s�hл�>���*�5\�Wb���ԧa�N",�w�;#�='�R��t����*�ZOW�0�.5ʷ��� ��-V_�f����Ry�$j(']gH���
�w<�C�����JQ��a���h�ع�{;����Y��g��to�	����r\���5�]�^�#�#����"J.J�ۦj ���B��r�����&f�16`�0Q���Pꏔ�Q