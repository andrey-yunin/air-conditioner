��/  �O�Ki�o�	(%�(�áS���R�?�$��1W���2Zpȏȁ��,ɒ�3a��p���VD�q
�g,��NX�mpS����.z���rT���Č�l,�J1�"\ʾwj��'�aV��5��g�y�װ}��1�y������ŌФ��δ_��ߩ�b�򰪋!^�0d��o߹���ɯyw:=G�`�9�PyCE��8%X�7	]�*����pogU��(~X� ��Vrv����P�Uh:l���V�	�$���p�2��_1y�ȯ�u� 4�D�M��hݿDI� 6�pn�l�!`' ��-1�=<H_6�n����rҨ�ҕcπ#L���)�yPk���l�5Y�.yIѯ9��6<���e
���-㘸�>4���)�O��K1,=^�h�ϡ�=@=h.�栜v6z�G,��6�� s|��~#7�gٯ�!z1$������U]�|�s�k��g\4�&���NC��PUm�u�^ϼ��0��C��w�f��!����a���}��7g;����U[���Z����R�{c9�wC�#�kf�WF$��qh��Pz&h
Z��
2��mw
�ʭjoO�֖���X	ɫ?hB����>��Ix���*^�W���8�)�d��������Ȩ�fO.H�����)��]���Ȳ�g�5���D5\��r�I�0t�8K��ز `auI�$Ӷ�n�r�m�k����v�o}�.�oN��|N��}x��gil��ί���Ea�T��CH�A�W��^[d�:2�!����A��Z3����R՗z�%Z6	y[3��#�P��}t1�v�]"���ڹĬc�_��Y�0ެ�z�͒<��Ө�T4�Uc��K	��fa�<����D�U	"I��w�oU���h�"Q��}q��Z�J�iH�[���ʂ�W}��h}������eb���� ���(�^S�i		B:����d����_ E�-ҷm�qn��dk���lA

nm�S�۳x;�����	6im���|�Ґ��͏?談�JJ��T�#��BT�1-G;�
���3��;(�C���BǶ��b?����Vy��z�ތ'�7�3�.L�B׶89��UB�ȟ�@�u���*�»[���<��4@KVLd��.}�1���u��"�J�g��˥h^�)1�
�;��ܥ��w�T-�!{��\�J/@G�a>��`������3L�6�2[��j����bEN`DR��
a)�Np�a?q\T�� �;=u` ����DY�l�z�q�!V7LslIת�}
U��X���w5�t�L?r��1�P;M�q:��E�o, ��<}�Rŋb�!����Z��/c��3���E�o�ZX+����l[�4�Z���� �$: ��*��5 ��ñٛ&9����6� ��_��	�?1��죫I�}�J�J���
��y�9��C�)�������T:�	y5S�w���� �������܇#8T��[�Ȣw��DZ���^�����Q Qag�h�
�`�Y�Ɖn�
��o�T ��^j)�5zDR
�Vnu �v��r� 7���\R9A�����2����@9`��)�j���2�r��:-,�G'�GO��6��{�	��O�m��,`�+u\��������ٲP��!*�[�]��SZ��H��pi�!>�魉4�uR#��EKXI8�^�z�s���rϢL�z#짱���94r�P���ÝC��Pe���7AW�晣Ĝ�p�G���z�=c*F��$���L�T1��|�h-�������s���>�H�-�s]a�$�����ӗ:o��������!�y���=h�HLg�|L��-j9�«������g7T/�4G+��W�!��%=`����<��� ���5��롔��-܏TDܤ�w���"��d�?_b�	���} �� ��(?W{�1Qp��#&���X��aoV�X���N�o�%(�Sf� ��	J�xf 5�FX�m����.�I��x9C@I^�V��aw2k����'sߙ2`���{u~d�v�X[C(�(��cT�|5��cq������L^���Z6	S�c`��Vgݡ� 'D6]x���D0�t�����(�M~nÆK�@�(ܖ9;�!#�A�>!*�}e�f� ��6q]Z�D+#���!��.e*1!�wQI�i�����#(.ZGY4��,�������<��ը��*������X���8٪ۛ����o�4�<~)��K��{!_�E�=gU �t���*�xaVZ�q��¨DU� ^���L�ކJ�/���d6�WJ�.���fB�K��} �����A�F��͋�;�����)�|fȓ�)
B*_����x37�xܱψ�>�ޜ+i�OVR39��
Z�幍J�M�Q�}��J�bwZX�Rll�0C�k�Lj�W��
S�E���NV$PO�|Z�-���C�t4���K:k��Yd8�+��)�Ih�i�MtX�w�A�M����.^�'��KM�s��b�d��v&��'E���ӏ��'6�l�L��;m���=$T�2 ���YX��m�뗹qU*�ΥF9\{��R��&y���I:�T��5,m�V� �26 (0*�'EO5��RJ�� ��%��$~z{����Dk%��3�I�{�.�j���;��r��5��H �k=�w{]I=��f_�UAљ�]�D/��ⷷ1�י���Ԣ�Ijl�	̖������{o��)VI���N9V,��H�m�҅��͐�P�Ƚ��J�Md���q�Z���]?�sIr���ܵ~z�����-�̓��=W��Y�%���O�r�}��J����:CAi����@�,�9��9�-�wn�����~�8n|J[��|�W����,A�Mp5�5>0�U[ ]r:Ұ�
k��wQ�LtT���y*��/��N �ʸ<Ԇ��K�\!ڭI)�b^�������@⾹�=��ע�@Ī�e>�=I��A���3����y���V��작<';5 ҖK����A.��T"�cG[r�j����*'*�W!�r"���d�����v]���=�0��CM�.t����qe��^�zj��W�~���'S5�	I �%�J_�ēJe�J��q{���*�m<7 �Q��Vc��Α�Ş��$52�
|1��QJ�4�A��t�Tck��O�<f��	�ᗚ�A�/K������N ����e� w�<}�w�(r|��k3�lħ�ʛBB���"?�A�@CR�X�w��|�nw��;� J��\ �46���ל��4ټ��z�X�폾�1QB&Dߺ�E�&�mm.OB�z��V���b'>�����傥T����C��g�K-���<5&�/�K�|bM�NQ|�*�֪>�;}�ȞB��Oz�Es:ib��,~ڕ��^�5�����מ��ވ;L|;5��ǫ�T�#�aW�L���j͙%���hv�!���X�{�ek�b�G��
��z�=��ca	t2J˜����_X����;�"�ʕe�2����j�<�z�CW1�e�~9w��b��\/y�J"��&M(�@_j���Z�b����E�/1^y���u��1�n[7�^���9]ox�pLsȒ�Æ����=��,�)�:8W�ĤXPL���2�eq�B��yX+��#�����̟-{T!;)�V���(n6:�s?��2��X��7=�.w�N�;U�'9l�8�(�`��5�ۄ+o!��fM�c� ��ۥ���"�}�{�]F����;���h:z_4�;��1M�O�ׅ����Y7�%��s�zMa���=����:��]�aCN�P<3���+�<՝�������\#�Zl���UƄU�J.��B4dp�L#��H��}�M�Hπ�9�x�gJ���to�Z�©�X�p��9IA+��������e�D��J1�7mE���ؖ��{�?C�J�=���X�i��"m,! �k�B$�i �ҷN���}�x��P�!C�G��˱���aB���{�͌(2��Jf3��K}���ʀb���8����I.k=�ZQ�m�b~�{B�Ϟ��1�r�u�5��~�����?�<�o2+Q(ء�=A����bN�ɩ�!r D!$����_�@�����	S:1���T&�s@��:�o�<�]��h�H%�46xz��US�
���&dn��鶏�,�}����Ks=���v�mد-�=�f3&���r�N�$��߬�>�Ys�I�u��9�J���"ʛ^�D>߳�ohoPglU�o������Z�Y���ų��o���3틅����J�A���L|�mo:�>8���t��G*��W��Z�4_�#�K)(�Ť�J� D��
}o7� �O�t�ӰSP�����D�.ؗ����׈��4�
�E�Q�C���g�˿IM�0��ɥ�+�%�a��]H5\���DT��� *H�M�J9A������Fd��I�|��ϗAE;yjQ�Ij�e�{m8��SS8�0TD������AT 	'� 5�iE�ÑGwGfc���3?�D[:�&�4�`��H~SH�A����(����Y�r6	~���pv~��TՎ$� �������v�VHt��* �L$��V.?:*�UY⃌=����S���20�A��cf�j3����~�L����l�x�!���ɓ#7o�3�,t��8���I@ʷ�����NJ��=�V������h�`��r�@U�/Z��VX�b�p呧=��z����5���n�K�|���EV-z�C�!��R��G��~T�2j0K� �����1'�"N�KIbo[-j2�i��(xW��u���	\Eg�X;b9�=�[�;	��>�@���1������U6UӋ��l�y��kf�.��ۚ����)��t��9U�I����8��	���U�[�߇�\���E�0q�.|ڂhӻM�0iSR�ʌ�ߕG��|�Y���� !�/���E���X&��K��"�Vw�IQ��/�T�piQ�9����e縄��9
6���|K�Z\�h�Dy��|y@��J� g�}���lD3����q��e�M&N�1h;���-� �S���tU�a��U�(�,@G���\�i�wDk3!	�E�P�{0��FD�$��uHt+�4�ۆbMQ�;i��xΝlԲ�[A�)W�;맾,8WD�� $��WgܖZ��'e�)��g�]T��g�2�` ��߷!��{����6d���6�_q�#���`Q7���B��<�$
�fX]�:KS�8�iv�^���,�T/�JN_�x�_�<[g'�(�疬�,vz<2ܡ	����&F�NZ�y����ϽD�&��08-��"(���m�����on7*�(��ćs��t�&Ԟo��1_���Cu*���7P��fJ��� Hu�E�v�|= �t�ZqЖȹ�Q�I���/��>b�Dv��c���w��|�H�߭���j?����MAt{��Չ�*ӭ�yKm��!��	A�����#j�k�H=�S����u�F�+�IUnD���{: n;Xp>����ʍ�
EX���G�#-ٳ^`��:���������F������NmբK^T�`�C��vV�����NC����`N۹h��>(l�<H��l�ii���Ӫ��Ch1�/\���w����jz�g%��%�aGD1F��Z����-{*45����o]x;> ���wZ��JR�X�m�^=P����y ��g��U:�v,��f��|crrw�˲@���)��,���$�ht���"t9x�����U�@~d�~:�ࡕ4Բ��� f0L�
<� ٪���:��9����2����t�^���3R�H���oI��r�ف�����,���ߝk�@1�tT�F����Pn]r����꡵�hV�改N��^��4��ر����߰(n~�0v��t~h�,���lO� 'j��,a�'��f�"eb���\ L��z��=-���	���}���ۡyS㌁�kZ��,8kd��\<�#I��o(@f���yh�;s��'�n��λ�+��i.U~�d�����V(>?V;L�#�&6�1����9���HZ�=��r7��<�ѳ>��9�qʜ.�(���F�i�Q�D���zY܅G����X4(�o�`�v��[�5J����턢.1Ӈ�6	;l[��6�Le�i�[�K�(�~�Fv~5.#����y]ıDw�=�s��glƯ1S�*���x�k�>@��y� yi/JI�~>�����Y��I�"��{�~���C^��ײ���RA[IK6�3�mZg�ї��@�'5��)pRG���f��@���*t/���Ld�6}��~,�^l��b�)짯c�!��8��(�56�gax�͡��}�x},}�}���Gb(@m�[u`̐��N�5Ga���D����]h�
���,*�q��ud�H�V8�\ުq���b��W?N�����r��,��RP�NܨEy§PY<�ȭ���m|�e�=>�0q� �x�P�����珥G��QJ��*Y�/�vb*I�߀3���bE8��	��9�lj�$1w�_t�1�/f<��E��CZY:d��6$lǵ�Y戩_���|�IH�}�ᶐ�0Ċ4�X��IJ\���(�T�hYXk���*�o�9���4eDC\tbBV!��);h9b~���-�]���?u��B�\%0F]��d�j&�X�����ظ��N� C%nP��-�&"�%�Ǿ���F'V�9��žD�ͮ���؁�4Ϸc�W<����s.��
�ܗ�$z�s�K����ԭ���O���@4�/�0�nO$q�ǋ�a�*����)�v�����C�1��:m2�/��qQYe��yCK]�L):O�����0!��M���]��x-�yO������:�Xɲ��NR�7&y�x][aI	tɸ�j!���#�io�Rʪ��	�ކc�PP��(_�|�̖Q�͇�l؆1k��I'G��{����1�+V7:n����  f���`�����w,�� ����V��bBs�˒s����NU6�U�1��]�)��q���h��f:�I�m���۩<Ь1�dY�Ia�S�z�?�6��	^��W%�w�ڏ��ac�L]����u�V�}$J�'��Hz�N�/K��#�9:�͂�!z
2���{<ۤ;��k��=�1�l9?@���V��3?zѺ����n���<W�X���~������h�x� `���m.N%v�I�$
N���#|QV�bS��@�ZZ�O�7C<��ݴdo�<T������i���S�:OKL�����*$y#��П�R��L:���h�	���t����n���%9���^攛�6�o!d�����2Ǵ��	쉾�����<!1�o���N.jw����G�W≙��/*&ѓ;6��Ҥ�Q@�Pn2�BπB#�d|/���ο���'��	Z����C50q��1+��ȪiS��F�-�QG`?�2��Z"a�=@ZQLZg8m4Z�+��^��(��k�6iHYfP7�0<��L�����埊	LG��^���mк�Et�R=1J]Ry?��
�S��^��
�h؁n�D����K��c��
� �E󨍻��w%?�?����D�UL�v���ο�,ք�.��A��Zߍ���P��H����
$y8�էt������D�a�ˠt�<(|f�z#Q��01kD���z�VU5����M�b�K��sܞp~t���ůUFd�!h�˞�d�;���q��Γ.u�x���-���Ŭ�D]������=��h\�ԪCqFƙ����P��m��\�TM%rD�ڙ��|���>���w���x{�SS�{e�	�k%+�C�����QUd��t���'�4����z"`��m�,k1g|�ǮG��L���Q�� ��	��p�/d�|.�"� �=J&�W�U���nZ�q�Y��ƱJ2��Q{Ԑ��2A�1�s)��_�ҷo8B�C���;)�3��<EOGI�z����U~ȄiF�BA�骙�5���GO�F-(�б��������Ӕp,EIH��UTi�[�o�"����5��)�n��..4�p\W��'P�����r5��o������Q�����ђ�E���ο�J3`�����J[.��E�����(����?��9'����%HE���05�L����Yi#j�?�ٲ�~�5��|_8z1A�.(��Vգcv�?V `�N
��r��"g�K��V�����@	x�l��
�b�����Ĵ/b{���iGB�c����	A�sF��,�n����s`�klg���+���dC�N����t��<b��w0d�!�J��N������A�.d��n�@�;�ϓ�
}��2轎�\U El�G�A�9Vq��x5���~��W��R�V�Jd���vu����j9%�=��:/����E��<�E���x��wT@��2Ly]O��2����zA�rQ;���OC���g5:�SJ���6�kA���c�W�)�!馩�$0�0�ߨ��	�jU������4�{(�$!xMq�`g�%4�~�}�����$'߻��k ���Q���=�d��H@���+���\��]�P!�g_�d��|��N�� g���3!ӲX�MZ']G]�m���`>�j��o>2��ܽ��M����'�gԦ=����l��\R@�����.@�-Ru�~����Ԓf�(a���?& W��:wr��wZ���s�5{�<~�Ϋ�I�L�ܤ�
�b�@+�a�̣�
�a�Q�o�}~2�������W%�,;[���3=��o����ow��
B���_ql��n�0�t�y3oS0��X�*��\%ǧ������Z:ۧ�u6]��d[����[��/�8��	k�����NV';,KP��F_WL��-�p��v�V1�5�U򅓧bϱ�_�k"�{@����N���5�@V�!�h'i�������Mh���S��[h�t|aρ�6�j�z`G�:����j�Es��p4��^�F�VR�y��VE��g�@��)/�ί���`�~wP�o���$R�r�`"g�w���y������ÄW����°V+�AE��?��ÍM��3#���Vȟ���vlH�Ƴ�֏/�b���v�
��#�%�*�A����e�+�JB�\�-��-j��i�%Ur�)�hȏg3zx��#rWW��i������Q�݄ɾ��.yO�]��u��ca0��1����ݷ|�vx��G}	�[�2᳛�ӣ.�6�"����YV����΀w6�����OC����0f͚�W�wE���As�$�F+�D/����(Q��P�x�m^�R�F��՝]�z]o��P�w?���\��!�-i��{\Z{�� ��u	U��@:K�.��w�2��t��������;"����u�^�-�k	�}fD�]Ș�Eœ�	U��k�[CAʯ_t�X��ł0����q�x��G���9�G8�4euSJ}P�����\�`�7��Cs34Ym��Sg���1����6k<����#�$YQq8��;@yG~糝7���4��Q���X���-��.]fY}#pMȤv\D_
}�-C���+X�K�s��;�k��{����C����4ΐ$T�'���p�r�odA��d�yܭ{A���^oyz�8%9�,!\qgrPs�u@��@��7N���錱���K��I@h�'Y��M�
e����=T��x.�z]�8���*����x�"�b�C�i�<�U�5_nD����}��r$�KW|>��̞�|kŚ�B�?ek�)���r��MÒn��ί��,)�S��U������u��>v�>hh�b��aɇ����#�� K���s��y^������at�n&aX�%ҩ��<�}%�M.
�?d[H�2�4=���j��"�����եٞˋҾ�J���Tt��n�Y1�%��='�?y�c��]�����%�LĖwtB�Rй gξY��Mc�a����<N�q�w�<��Hζeܾ�*nI�-�keL���89�0�Ԣ��))t�mkz� }�Ť<(V�KJ̕�<40噞ׂ�	����U��F��/�/��G�`�t`Ȧw@)_nv�U�[��9�,�+�����&�d潐��x�X����u"�_T��(�����©��n�=�qI��뗏�]0�[�a[��T�Ê�W�˼~��w��%ɵB�l3��<V����'������D҈�z��\�R܃_$o���}�k�Q������o��M�,[��a��Fު�_Ӗ&RDezD�۬�0���${�GT�e��|Hk����-s�����<V��BR1p���`8#���e���>w��1k_���җ狇���� �Za��.����j%�	�'�x|�3���D���6T�6�*���PM+oYM�/�G"V|F���N8
^v8����3�;�R�x=`�s�*7QOv��q� ��o\C����3�V�@N72y��o���MG����m���o�ͺ��ue{�|��΀	���ǅ����i�sv�%��@Y��ߊ��(��R����Vul�V�<b�A=7�.�J�������=�(���pJv��Pᅆ�Ha�M�{
������!7bQ�}W�·
�M+���zu{]w�s�;���N��H�9�l4�֤;���kJ��j�J��{�aZEr��D½	�T�kgX#�z�H:���bĿ��kP�%�n5�tx�K@���C���"(!����9�P!���0&�,}�3�x�	p���B��;�,��� �w>������g��DN����:��n��n�=�����^�6Z���,-���Y��!���D��ڢ�]��FK]���:��(���kL.���aa�\��$j��)P��2�:���l{wӳAHYt��,a��WT
�� yaN��!�-��<�6MJ�7�m���>�hx�5�,�*���ॆ<�-�Z~�O}?EM��ld�,5*�zs詩�Jk(�v�ʾt*�C����B��	� 9.�I��2��S�[�d ��T~L�h�z䕛(ǣ����ᬞ����
�u�%��Zu�k�w��L��\&��Q߿ŧd�_�pDEgȺ_ށ�Y�������zd�HY���F��ӳ�6	`CY���g>�T#g�!��^�h��ݴd�o�Gɽuq+@¶�p���>��Q��cu�ӚCX�^�V��x��3�q�ދ_$���q�W̬]��윝��P�\�9���_��g<Z��Z��B�38@?�e)�vu�UJ,\�3 ��fD����
�k��p�{Ŀe�Э��H��V�]��M���7�im�K��x~���y+D�-�¤m�f�v�C��"f(�;b�~��&?�/��=�i�&m_�JCՍ��b�k��n�0�-��� ��q��������s��!����y���2�6Ň}�B�O�gz-PVR��~feN?E�ac��-`�2���o߾l۴��F�����X��I|��I{�#��m~�������i)���
�;��U�Vj�0�D���l�ip?��V�RB�P>�G��k��s~���!Vf* ʓ�u!��1��Tq\  ÃY�}9K�9!�������\�d�s$��fK@��F����B
�Ap��s���w�qWt΅+�KU p%��˒��H���e���q�}~�l��3�N$��M��ҙ��x�/(��+%"�ȪcU�R�u�?�Ǝ�O�BkC��6�G�?Ym��J 1�6�1o,�*�NU�����PW"���<}UCp(�V�����
ȡhBF�Y�KG9$�M���M�ڿ�߀�0��-R�"��7��J���k�/R�*�X�θL���9��B���R�3Y��
nSac�|��؀��+W!�N���0�g0:-OE��Н�U�4�d|{(��"OuygwU$7|�Я���F�(zw��Q$0���`�������C�=m� ��BC��/��P�UI�[O��Jfoz��=�$�$c�jNO#����;���2Qpm�wDl尜\�2W��>m>��o6e�
���".O��E [ϒ�cyH~��f#�i���{�C*��&&��ہ�n[b�8�԰�H���	Y��å�Pl�v@/N*���:p2����E�ؑK�B�`|@R�G��^�r��)Y�����D� ��<��&]Tc��������H����s���"��n�������d&a�շ��2���N�,��B�4���V�MҢ�o׸FbKU�*D�0��NR�l���r��hh\
����q5s��	BV0m�]��v/��W�����9��f򕧢�cH�+J��\������6�g8�:{�5���u4��x]��ɾ�|B�ԕ}�YnB֋B���J�H�kJ�DQJ�F�ǆ�������8�3`�����d{��C�Ls�QC�H#]�w���ǁ^�wo��Z�AV��{q��Sn� �����q]�H;$�iB�����`尺�Z���p/Mu�<5���n����Z�]�}��;C��uN��5�l8J�%Dd���B���˘��������q��f�[��~�ϊԀ��Lz��H�D[G�զ�a:�SV��@�Ix Ns ��kmό�k{!���1t�]˟���D����-r���[S�.��Sv��/տ�N{���$t��:�>���E�ty	���pJ&��N�k�&B>1k��}.�ʬZr��X���oɭ\;�}kQ�H6"Dcۅ\Y�4I��j��f49w3^�n*�5:�Q|���6�w�t��z^���u~�/r�<hC��B�{"W�5��P���9�֫��m#���y�͓$��g)����3�"��ӌ�u#��B/X�~ֽ��έ]�ߝEtZL�����U᤟bI0��@@�8��|�e-�_� "�\0��j�yŧ!Y��b��Z���S�3x��o<x�5���D<F�R�����At9�P&V�6m��V��p��gv4B���?��/ #XT�BraX�8��m3wpW��b����]aXh�)����;�����g��cS%�t���uB\��DQe$����2jO�"����m�4 �Uj�D�}��!3�(�#�*��7St��D�h�:��ś^�r�j���Iꊚh�!_[�}��UX�G�:����/��|%����s/" #�m����W��b���}f�6��+�:�V[���~5���0�����A{�wn�Ǘ������)�$����4پ,j��f���s3�0�<��]pJ�`K�����\�`��t�� J����(}>sQ�������ٖ�k�V�!M�*;<�.B��fb ��ӑ��ы0+�&�s����jv��l,�p�oQC��G<<\��jS�P�	"`:���D�#:�j��A����_�1����h5��
��0��I$6������P�`���%R\�L�x�Z��S�cf�}��o�bf2��c�z��o�L� ����K�_�-3Ngw�t[J�a����jL��;�v��'q�bV-����Za��m#�(��ʥ�ls!h���[�u_�UL��f��#�K���8�$���[A�w$n�q�U2ڷ��������ZpW^n�͌��}�>1�.%�{�st�?ֱd*��m���FK)�b�~�3*�jg��Ma���p�+��w����2��C�w�ťX����1/���$Qԙ�ފB��0�Ч��i�܁5��x,i˽�m��!3�P�3���W��P^��f��̯�%���ipWE�`�->�R�
�n�HC�O�������h�(����&��\��&��^�QG�qg�\���X7D�I�䩢؝h5���G���`�퐍��*)Q���AB_T�-�E��&)D�ɅE�jԉ�&�p��5"�� K��<�)!^H?>{,���g�ɼ8h���ǰ�m�]k���j�|��͌��}ǂ��#<��]�ת[JO��龯h򂟹�>U5�W��v|�E&��nƠ[����!����\��&�ɤ�q���gLW��i	����P� ���jm�ъ�i���1��Y�2wv4uk�A��rt�?��VdL��gƳ@�Wс�(����g�x����Nj.v� �%)��D�}���/J��P>}5�"��uA�z��3���(_w�+j��6��#6N��Xg s��ZV��Z�ǡ���`R�F��x��牸��@l�(ɂ�ܪ<�����.�50@:���6~.U��
S�٧�S�)�h���da������5�@יg�R@E�72"sMSv�2>���Β�>i��W��� .�=u��EU6�*���Z�d�Q��U4�7���;Fm��Y�Fx���-���>O@m'�I���0(��}�c�(���_�������7����_��!�D3j�0���2�g����ʁ���֮��a�|�����Pj�T+�(��`������
��2@�"������Oҩ|V����x��w�K���/a���É��a�6��d��_8�w����=~2)��4��{������ߪV�{���-�6t�K]N��5�(�;	~�@3�N�:,D�2���gԉ����S����>�0���A��[Q'��/���&�����˜�t��,[^�{�2T�6ޟ�	E f�����~O@⧨kP��c����HD�(�Z_y@,L��#S�^�֡ݫtt%<�l$YU(<����ߓY�8�Kr��ﹸ6���`�{��RF�d��=eX7&��T��ԟ޾
��3T�c�����Q76s�h�W�\���8� �:�Y�S�;�!"��oy0kIK!�V��b�z8�c4o�Q�{��ҍZ�[<j}���ִT�lE@/�,��k�����2�306e(�4��D�׬���`�]���P�Wf MHa�����0���x�$�<��c�yo�J|#p���k@$� ۈn����ӕ�	a���[���Xh2���@� y�t9Ň��Y�Wen%��ل�0d�;
�s�$���2��0���2��G-��3B"p���%e�.m�S��Gd�K�����ʞ��	�z�[���,��O���M��=�Y�{�VS_��5�cx�5�����D/�s��1\ՙ�&��۽-ū?5y���H{I�dN������:�J�M}k9���j��k�������z:���UO/���j�o����\��FV-#� ��ܾ8�1�<��CWpᰉ��[%��o�vg�?K
YI(߀,�EI0��}5[�5>���Ca#JS{+�~q����;�y�T�l�9����s�՟X\�	�wL�������5v]��8հB�ї��Yo>��'�����<����9@�߰Z��y�٭��4���/�_�t��Ɗs$�@�|��,�~w�u�P{+ܷ;�v;%?����y���~q��t���c��V�F">q��%��hλ�c���swyd[i���f��,��R�=�y����:S�>O�+��q����w7�ȫ�9���҄[k6W���m�:Bӥ��w��� ƚa�ஓ�nI�B�Q�ʭU�Q�e%��<E��F�z>�Ӱ/���OG0�k����������Yڈ�g�4�ETG$7���풑�^���q�������9�ʼIS,1*�9�>�@��7�k�XWl̄�TV����!@���tR&"����#��`�K��[*/�<�Z؄�fJ�$.VVxb��W��O�K�5� ��$�jP�'�����s��sU�S�d�=�s�P�a�&� c�#�e����H��E"w�:I@��U��U�xU��1�)��鲂���Qnx�G����g��im�w�&�5I�W�?���-R��G��=q�s5nd�0隡IHW'��re��� wn��k(�Tx�R��ù�R��)Cv�����F��)�4����K84�(\g��&>�}�����Yr�����f$�ό��p�����qV��� }B&����X9��J��=�yK���uC�(Ss^��܍!#��c\���=ٟ�!q�Ԙ�XJ�Ü��/S8�x�2	���8�}p�{��\Vψ�i	�� �:I�!Ʋ� <[��eI���s�(���=ͬЂ�����?@E�go0ЉI�]�*�/O^�$��}ꙝ��Z�(UX�y�\�s*OP7�]9Y)��?�ɯ�/�c��V�u��S߷I��xse.�?(q(��OZ���+_�E����Oo:(��m���o�������'0Ĩ���:	�f=".�}{lWi��ߕl�=�'���8Ln:���U( &��k�P�zݑ0yw-�`C���p�й22��{<��p����s�x�4�b��!@6;pÇ9�;)`!�O�h�[%�D(�x�Wo��.P1
��˪�F��v���j��J�q��6R� F����oə�So5+�T�8cA��9BB6�g��%dL!�J�|�`9vJs�d��P1_��ms���w��9�s�����N ���Y���?�9������~�Fe�iF���'���`7�@
���I�w�D��D�¡��j0��S@���0=y���m���xBҘ�%���=GS�&�����z�#T���@�y6�������T�G�!5o�_���M�|u��ٔ�)LO0�X�wQ����*���7Bn��&J���V��-����|%+^̅*�0Hu)��rG�s�Y���p-��0�����w5�ޏ�7A3�Hw���ڸ�(M�=��b|��X�43��,�yGM su��0-s)�����lZ�M*���i4�)����˿�t���6��s�?G�I� �,7�Q	p5�:pI������W�6�K�2����
.��5Z�F��z�����[D�z�|�`N����zA�0�Q����Ǩ����Q)�*}�.�cD)j��cpA��qc��h�!��hx�Zw�Uz*�wMJ��\_�&Uހ��S� @�8��f uؒi�u}��;-�	
����H����9. �W��(+�a
�t2Ά�Dp[�%���roE�����Y��������h�Y9uQͽLL��&rp]��7V{�{+wN�[=���X��&7�L�C.`FM����s��b� *m��`�sg�U�!ms���H�'���'��LD�TA�_��2u�}��Y(�Bd�X��e�V�̚��@(+�{K&4g��[!������� �rltAc�K]G5ˢ����#xw��������=	�yM�����x1��݈Ll�F�ץ�3a'�㘂g#d��������x�!]�!xm]Ɲ�w�t��?S��jl(��bB<@+��O~�x��v��W��H{-�d��ԫ�={[�@Q���eIqc{�	�d|��z6�*	P�33�cz��z�p�]�"˧���Ta/�e1�W>4���]|�ظt-��7p֍�d'� �8�J��a}*�ڥ8��\
�����]��S1j'!�ϯ]�2�i�+� �q:Y�� Q#O�X��&JP�^����x�w79��;���8zY�[�L:I�˭߃�O2�,ǀh�s��3�[�L�bx��Lt�v�͉��	�q=Xp>�蠖���\�6��%�"����*��0#^��Y
��O���)"�8N��V�j	�X4D/S�N�~���pŦ6*y�>r�L)&
��u�+�c2;d*�Jv`��l�~&�ؗ�����4,��3����G�#�.$�U�D�cp~�= �=6Җb�F3���r�;����]�M�[�q"��&b�q|�ɯS�d4��}�O�&0����mg�Kn����O�7 &ǩ�|L���i�Y�y��+04�%��Q�$V���#$���Λ�����!�;���D�Q�YYh��������`�g$�Zۻ�%^�G1p	�r� �ޒx�%� �q�{�� c���Ī���81P��v��Re'���z�SY��?����G�ESFZ��`8�������o�$��Z���=�_���=�ޗ#���k:�D�C�1���"�="���&����$�$X�)���-��	�7U�[���O�
�&�S�Y�+h�O��s�=łJ��-�!<��=׆�a�<�U�07��&�4e^�W�o����N��{S��  �I���xY% �ݼ��͙{Xˌ�����ps-����P�N�K~�Ǵad��r`6�$u�]H���/u-`�<O��d&Kk7�a]���t}�L���;9:��r�ʲû�׻�3��B�g��zp},�۵moi	0�R��5�n7y�KN'����R|�[���1(�s�\�|��	p0ڣ͝y���|,�������9~��Ҥ���n��O (�:�Õ��'f�����āJ$qunh��a�,C��\�r�jV�'c��!_ݦ�9�ojo�m[���ǈ���z�7]R��Y]�=��꟎�p,XK�JW�.��8��r`���(��ԡ���X������^�-:��44��O�|Q�Й2�d3�����OV\�P�4u^#c�xM|�}�fm�[�p$�3-��-{�2�����`ik�� �C��Kv4�b׵�c[9�M��g��zK�V!�m�K�PIRO��z�m��+�Kؕ.%�� ��4�����{��+�=��o5����>����X����7���}Jab�aA<��L>^jVt��tĞ���UԱ��姸YQ�Kjɀ_R�>\�oA�(�eR���
��m�L^����������z-�����L�k4敘�����h}�կ1�ъ��~^!q�E�қe��Bn� -q���hҞ ��������t.> (�|���VOU�E�{�=N{O����{��XG�s�~D�Ch���(?(�3��n��h1��6}�6�\�░�+��m87>{u����e�+��8jSU�>�#%5��|#P��� ��؉�Z�b �� �0�c<*��D/K��|a�שl����O6�\c�[p4fq>�GZ� ��?���j���sY�`�����4�4�V](�iH΋��R��WK�]�ؖ��͒l��t��%�_�HLvz1y�H�P�мP�37&���ج�Z�����}��zz�kU�=���L�28�鼢W�캃/1���D'����ϣ��4�H����񜩈|�-�O|r�ӀJ�_Y<.��R�ĺ�R���g�:�O��Z��J�k�|�S�i���e���L��427�n��mw�j�
���&YX0H$��ft�y�ò#��4�1��I��6�t�%��i��KE/\Dl��9��O�~\�	�a�6�P�.�`xe3]�����H}�ZF�W�0IK�F�36Qƫ���y�Z��W.	g�,@��3�x�\h�a�QT�D�%)���,�m��kt� �j8j�� 5���S;7���G1��1�A��w��W�Q5�Ѱ���D��o)��������ݶ{�$B?�~�����w���x�ꫂn� ڠ=�� v���q��8޽���8��E¾-�1tc;IU��E� ���4��m�$sYk2\	0��fH$�T(���Nf2��R�-�B���J���>gj�̻�zd.
�y�ѣ�gF1�Hl�yȼ������PQ������=Y]]+���`�l3e~C��~���7������YA~L,�SԧC5�Gr�]LhOZ��U������=]�[��\yV|v���=�Q0��lf@ �)�����u�S�ښ�P_5(�̺�9��f�?Ϲ�/�E���o��nCҶ��3��*SZ�߹�T������/��Y<�7�-�'�t�W���V�3McN���h�y�վlW_����]؆��T����J