��/  ۷bꧽ+�m{D��:���\��-&�$���[���6������������3:Ź�iukqZ&ݔ��D�T��^�`�n��9*P�<�u��x܎��9�79$>(�לC��G̎���o��+���g1�I=�R���q�<��آU��V�wDi;~���'�ǰ��!^�0d��o߹���ɯyw:=G�`�9�PyCE��8%X�7	]�*����pogU��(~X� ��Vrv����P�Uh:l���V�	�$���p�2��_1y�ȯ�u� 4�D�M��hݿDI� 6�pn�l�!`' ��-1�=<H_6�n����x�����dǅp��U���$�qɴ�b�6��|����0U�e���>7�/��(L�dՙ䆲�e��v�>ǎ ��uZq0��t�L�U�ϹZ�`�V�:C���hN�H��_�j��PЗ�����"s�=��� ����	a�8���<9Eň��[.����;�b]ēݭ����j��>z-g�@������@�e��Ѭ�.r�u�N��T��ۓ�6�������0��K���ح�U�Q�.è	��]B�J�|����w3��e+c9�Z%��v���=@��cn��5$�Y����_a�kE|L�tW�1hv���{��'8�9�K���'6�Ϥ��	h����(܋C��J���$�D�-#�We���{s�����l/��3P�2R����^
�q���v6\s#�ܲ��5\���S��R���b����u�Ot;چ�N�$��X>:����L`g�qf7&�ɨUo�-����h|��HM���P��&v�6���؜7XP��#�������������Wی�S��O�O���N��%�t$���Q�t���f!��>�A�%��!"�m*z�
 (O���1J��Վ� ��g�5�0��ni��e��a�s��+��C�����0���d���./�0B���p�bQaL����}G�b(�s��Ay�^�~`�g2��t5hC�W2�Q~sB���m����ÐH-��W�S:��;}C��3Ȥa�1+#�ټfrl��J�ٙ�b�Ӻ���?��j_��'�֋����}��j1�)��S=�z����П��h�W�l�7VN����EE�)�Mv��ב'���'P(�Aα:,���A���
�Y���0�jF��#$R�xH����u�$�쏁듴��yAu��tں�"���'�SA|�E5��Ƽ�N����{꬘�!D�6���9cy���ͨH7 �
o5R=� �:U��j�Z/S����Hj=��&k����w�!��Ӿ����(�5?�0ٗ��E�.'�Y����!Z��#4)��p� �J;������d[�<J�][�(��SK��ϑ�#�h�`/��	t�M%VȢ멣�d* ����(��V4�Λ�
�TG4��]ï!�Kwzzb��s��2?���Ť���	 e_mG �1��j,�n���Ӎ^�/�k�q(�{�803�k�S���>��F�5��-d��#(�ET ��HT�_��h�-V���I�f����~<p�a3&�F1C���_<����+ϡW��EI�%A�g��F�P�U,���ۻTW�qv6,_]WP��������j(LW�r(��_M$Z1�Z��v6쯘���'|p�0/c�]��$SG��1V����韯��-cOe�]&�-��[����H�B�s!3�z�jA?	�E�7��3�}����g�gZ��F��Ȥ3�3&����*/���+�Ȱ'g�P��U����ل��uQ��_�h���8'�#�a>ҝ�9e�9�qڠYnV�-�G�[��Pm��y.�A����-��z�'�j��u8I��:��j�Z4&{���Q����9���c$nP' �n��i�[q�L/PK��,�+p; n�6(����4�0�X+]In7v���״�}�M� �������������-��7F`c*�˯�E}�5Ǹ81:�#�ÖIhq�+^��/�����.�*��j����)�g������;4��F���g�8��N�����4�6�.o�r|��M���۴��ݛ��濡qݖ�
j`� �%�}�y�{��?=�H�M��-��S� /����P��Iz��KR����e�x�SͦOU���[	W�]6d�Z5�%��&}���w���8��ގu��N�o#}��Am�r��|��8�ɂ?���\��v)���#mq�iN�l)�&W�9��eaX�6|�L��B���K4�Vt�=-n2K�@�ܦ�W3�!�B6�V MY*.����uQ���B�(��Ð��0�߶,����z���ȜZVi
5�AĬ�C!Њ��9�ҏ�v	�5_��i_�����h5uw_�&��������G�ta��V��GM�A�����f9	�� ���vK�������X��F�LƯQ�3t��2Pۘt��MF�p����&R3��]5�;W=�ƒ�ii��K���z�Z<h�m?��t"jf��a�+=��g[�weqx�,��0�R�1�� 7kD�B��ౝ�>+�6���������X�o�ξ��N�]h�����$���������/����L���%5��L�x��#�e��);s֑kԊx�T����
,�����7��I�8��6�)�	�d�j���	-�r=���/*�(f���n3	���@���cj̯!ܩd��p.�mKI]_H�X�C��̟����R5��iN���A�5b�}��.�*V�Sm҈#R�O����;2��7y�x�{�xKVY���C5�]�����_P������w"r�x��j��P�슥��9��ҷ����T]`OK��SH5=̳,�gCVG�� �:ǌ�b�gwȡ�.�@l0���'�p�R'8�`��aI4 6eo���>�����bX(�H��~6�ty�D3>����s�h5�$��:��7�M����n��� *!f�&<k��q%f2�J���d	���/�1�k@9I�k�A�����(���%^x��м8j}�/��S��VoLS��Or���CZ�#"�v	���6�G��L�ݨ����(�D��rj�݋I/x�ݮ	��S��"$ey�[E	�}�2���gjܗ�C']Bg4�<���ڥ���KX���@K�(���F����V���]�,8M"��;����3M7TI0��#�Lg>��g��#��i(����0�&��z�\m.�k�U��Q�N�iʺ����tb���/C��$%���@z'4-墋�K�W��>�?� �B .�Ψ�V����&�"ai6	�9�|�z
�kl*���ea��Q�>�2P� f�S���6Oer���,g��J7��ۘ�7�(Q~*�f�
���Aٗ��},/ϩw�T`�\\���/Hp�[f��SL�($�{0{Z[~�+���vu����Z�u�DhԂ���.$�n�T���@�����d���lLBm�W�������2�6E�>������O�����;�J�sA��xWU�&�W]�M�0� �Wղ�=e�k�-� [K:���b���%�ة���L��x#�V�
Qb|�X�tX�u�	2�#� G�:�p(yA����а��҆�C�P�����v3��h��0F��6bۃ����R� �a��Y �����W\�¾[o�p�*>��ω�7�O|ɋc�j��%��M�lV��������
���IBxk����T��W� �8��<'AOH��Tæ���$���m>�XΌ����Nv�0��v#�CjɽT|u�ΔI )��KA ��&=�Bҧ�B���$�%5\V~��T�єOV�7�Ni�i�"�f.�@�R��􄐴��`Q|{��,���[Y�0z�,sBda)�a��(xg	!�d:mu�d�8ozۚw�����3�ݎ����$�|�y/Vb&ݶ�x.8�����!1��N죚Z����N�t�U�	
w���&W�{d��|�U���p�
�8��6��[HZ/�\���J��q6m1r�k'"�v�91-ۏ�G��#8�������vb=�^���L�spC,t��1H�&^0R��!�Lx��ǔME����U򏔭���h�����y��$�{:����J�����U���Q��<���e��V#Z׮�k8J��to8VB����G�1p�6�_;�av�T��F����H�KzCG���t���,��y�玛}��%t��&o>ޠ<1�%n�����u.]G�l���r8��y7K}Τ�g�y(� ,�ys��xˮ	�1�ؿ����,I=�����B�����P���ht���c/eL�D1,��%����b�$W5^u��s�;�'�A�9����A�p.�9�N��[[lR5'k�5-)!����l�m�H���'p�eW�bu��Ҹɚl�b��y���@,�vg�-�4�M��f���vl�K��v����*��G�����]2O�L+ �
����:�*�����+T��0�m &"e����@��p��8���"\�~��|ϙ�]e�9![d�~J$^��Nɽ��/U6oT0��W�
��c"��cL�̋���{���~�d�#�c�AǈE�޼28�7c]`J�l��8%e�����󃚌y �,P!��]�~�~�:"��h�c��vi�̽�ǈ��d: |���\a܏�g�܂�K���b�e��� ��m���O�f�XBR4��h�V�w.%)�꤫I�(^K3��*�怔�Oz����66.�م����rҼ��ιF��;�[G�43s��8� �D�>�_����*|n��!|!!1�7$��p�y��3)]>�D���5���Y�T�f��i]��	{>����W���6	[ f@�����d�b_j∘	rʰ���F���{���4$�1#���2���=��p|�����<�VA�\�^0nD�D+9�2e��405{�w��g�ɋtv��C�,+��fU�qOL������/w#��~,�A!C#G)�~���|���{,�r���I�W0��Kł������]���r�m��p'��'�ɬı���G��wN%�G�ì��h�Oއ��uE��1y(_�+�dI���M�z&AO��m�H�L��_�_Z��_��L���֕ڜ����i���q�;��CˁT�U��zb	>*�:� �ʿ5'�á6�$ܠ���J7@V����B�'�f��$���n��j�&�+��H.~j�����&c����8V�I��8骷��j&�/6��SJ�E!�y���x3�U�8��J����|�)�\�QP��6�Y쉱PW䙎�&�iEx9�֕%7!�%f�ęY���d+Ar�q����p��L����V��C��7��osw��ףUOѢ���P�Exsmn)�٪#�&S��%7�0�ځ�c0�Z�;��<Y�z�X}�U\����6}��բ�,Lk���;?��A��7D�h'�3�j8CC4}.M,�8����Ja$�2��	֑�yKhD���[Bv�5_duV k�Å�D�s�YfqK���"��%�-U.r.��N�j΍��v��b�s�k�h�.��D�a`O�J���SԾe$Hz�+�~x'��'&� w��� ?g|�^`��'\��m=(<P��S��s�g��.�73��v�c����'f�?a.5\x����*Z.�ak��ԭ���t�i!�c���|�y;�ʱS�� h^Գ��l�|��Y$|�0#�J�W)N�]~DF��$_f/|��ԹNG)3�����R�͔�ܫ����zZ �����;k,���n�𿄖��\9t��S"].��q+Mz��D�;����ʛ}��ʭ��Ed��r50&`�������u��"S��u7�#.s���[+�]��U��.
�]?W#"��G$�^֮2!��'#Q-��ۙQ�#�c+��V��n�Ġ�<���)��1rm3�>Y���9���÷�!��2�	y�z��:=��
�ɤ�������a��Z��p�E9��]�K��Z� �ߠ�"�:U�߾bE~.Hs��L:��T��.�%ǖ�M%��JQo�`�3��K�Z����eU�(�4^�Q�,��`1	���ux�]+Dⵕa+�Z�N��}f("��d]x��.����7Fj�ty��-&��\L��_��7W��,a�N��=I�`E&�ue
�x�u�]2��5�bp��"��陡`v$C�0����+?G���2�'JS����x��Q�)&Y�ӽ��g�4_�4C�~�#�_������Ya65��P�Cx���Cu���"�Α��XM͌���wqu�h�HW���L.�;%���@�������g�յ�u��5)�Hc(3�d]|kQeb�]`r���n�h's<�pm1������'�O�n�{�'�F�}���i�"j�w�L]c�^���*�n,kE�vE)Aʙ��v����oE�_�<������}#�z�Aeb0+b�����T�<�aaE:�>�|n�-
 aZ��mG՛��p��#�������U����\3T�5����LN%R!l����7�w�֛7^sI^�����J�豻��	���4�X���7��?�O�ͮVrp�Ct �"�ߜ"�UJ�nس!�Z; ��W���� �i)�ꍏ��z�fWDT�آ�EN�,���`��3djm�8�U!TǠq�3fx�I���qv�|$s�@�u���gm9�]���7'�)����e�ަ>�v<�dF�U����J
�G�ie%�ƂJ�0���OazC`qY8�t��!��fԮn�z�l�Ҭ��ދ���,0ϭ��/��hN	��%�>�F��6�F�KT@nT���P��r<���Z����}Jir���s.�`d�M���#�#r�h{�pƚ�,�R����]�U�	f���+Q�8�_���a�2{�4�蹸/�W!��a�E�گ,p�풉�����^�3�j���&M-�|�[�&=<�2B�� �GRip7�
K@i^~��J�#+%I{�~��5f�Ng�4~�mU-*���bƛ�32��p�����ͅ���V���9N��Iz{\{"{o6ѥ&��A��"l�S#��ʀ'�mo�L$��!"��}��J�s�E��Ugvi��gÆ1����B�B��@�J~�[E�ko8���+�"O��/͓��AX�z����(�y� �~y��b�~���T�ֿ��׀������^/��]��л���/3���[���giL������_зV&{}}��=�ђ4;��_h����bR���uY��y�s�H,���l��,�k��yA6Q:q(��j*|]�,�/z�_%���{�r�<�g\���g�tum����N�ڬc_!�>����v7c 0��JF�>>f��NCD���a��h��C*�a?����?3G����a�-��8�˃Q����S������4d�����,��2ԃb dW%� ���L�(���6,=�
X�ǧ