��/  ��*pҥ�6��Y-�#p�\K���,���V6j�ј=%��K"��Q���>���T�mW8���GL���Q����LB53`��ݰ:ޫ�>�oa3�Z�&MU�i��êR���:�P;�F��C����/o=˴�����jV�7��eV���+��~+α^��P7&����n5e�%!�p���B�\dX�z�xo�m7��,-D��fI�z,͢*2>P��RB،�$��tC�<o�����@6�R�2�| �`�y�y����>I�_Ť�2����2�Ԋ�Fp򞹱 3ǈ�qs��a:���'�z��t4x�8f�B�+�@�{�Ǭ����V3Cu��M3��! a���	�����_�J��r�4f��Fa}�����ΐ����᷷!j	Б|��D�6>�����5Ah�d�8Xe��\6�S����D��v��pT#	ր�M��b��O�Mo�M� ja_��G���i��C}�����8+�J�MeR��9y�矀(��ID������t�Sl����Ndݦ�0h��M��p�|��Id^��7����1^
�Q�J���C8��S����[�v���tX�<�\;�k�K���\��K����Q�X�F4E�=�xAԷC�ʔ=�k����g`���V'���D�8���:��b1��T_�t����I�?��}��M�t�.	��Z<��U���%(ָ��"m���e �ЕP�ks�.�CM
�ʚ'Kp��BcWн*��[�F����V�"���Vqi���v7��X�g�s�����7���~��T���:K5�	qb���H{�
�Z���>�o �H
HR��((���sd�q)�2}_����5MT3�Y[�U*Ꟃ���_Rk�^�8�dû��X9׎RT&�|n"��C�J*�~��j�?_�$�NY��#�T�Xh�j�H�/�>���I���Wj�Vy�4�r=�)e�S�L@��;��K�Ӛ��Z6˴�7Sj^���W�AX�56����z��]�+�e��^|@ρ�ٹM�M|I@]	����j� т6*���9� ��!����d-l��[qc�bH�b(�����!ɯ��6?�lD���n�A�e5ڿ��{��Q�8Ds�N)nu~h[%C�i�RA����]ĺ���>��0@��tu|��/Ԇ�yP�F�]9F+��xs�j�`� *���ig�?�r��g/�[gݰ��`{�5@��\���Y����}EϹ�5�����������R�J��e�乻i���v�e�]Q	�@o 0k�m͹��*-2��z�ɂ�0b;�$��*͋��z�:��g�X�0��!ȳ O�z���&n�(�*yqxQ�t��+E[�����F)MA��C!_C�f<
6(�7�`��k�&�1M�9f�N�6�3���V��N�0�\Rn<���R�C��e�����y.�w1a�����yU�˼����ԟyB��wT{.�I�ܢ����M)���Em4�nM�*�jNN[���'�]�k��Ĝ�6+4���i�̱��Ł"^2E�ݾ_�q7h�ة,\`�$�k�Pާ罚�U8̷�hLI�v94X�UA`�ez��,^�����>D�F<u�3p��Yz�]D�I�m��Lƴ�/�`���NpL��cYwz�m�mk�ܠ�}���;�f����27��RAU6*�g곻]����(�W�E����J�~i_
DF��xO���V��1�*͏�Hh*Lǟ�,�u��U�NGU7	s�G�~�=��fb��h��ndQ�ԬR..�F{��F���?��ܝ|�Z�q�h�A������ڷS��z������ u�%�qv9?qR*}+Knk��zܩ��Ǝ�OYvy$p':�Z ����ɰDO`���Ű�3�?����|�3�$Ǻ���#�����h#չ�l��M��'�� �r�X ����JG7�׏*�FM�B������=�e�<�3��F�#"_7Dd_x^|8(@�����nr����kpA�T�w�+��\�~*��P�e��gהJAC�� �[�e�)qܲ�-!�b�i�(8v&p'.�)L��,cF��Ιr��ǜY۽��،���BkX*02ʊ}�V��S��n�>�rv ��{�i�M/�,�I��˻�9�xwV(w�I�V�I����C���C(P]3a}������q�a^:D��V�]�f �)��`p����%�;� ���Iӆ�Z.��W $T�Y�u��������p.x�}�]؞1pK�6>�t�ZŴ�|y��-�K����Ѻ��P�41!�������?�WM%o"����D�03�(�R�E����"�)n���ޞ:��JZ�,; l�u�}�Í+*��]DM���w�G�������i�̨b�l�VfISQעR���8�""j3�&�����'q!��k}'�1L�j�*C4&��U.���;e��;
�]on'z^���V�G/���@O]Ġ��X?y�w��Y�
�|gF����k'Ɇ�I��K��BnmAB�H�WBL&���q5K�h��8i|^�����Ƈ��v�0~s�ͪ�
Z_��D1i�^ˇ��*&�B�GT�Bt�T!T��j���g�Uэ��#����(T�
�|hM�(��ru��g���ޤ4Q6����x-4e�+���#ԃ�����ù�� �nj17\�cTq�ϛp�G�)�Zy���lCr���@]{h@'��	��J��r�(����%�#~��3����Ȟ��,TC�Kɰ(�d�إn����u���o�����'�_ʁHwH0����� %��Z(��Rs���(��е>�r�!~��tx�5}~�햲!Q8�mLޭX�Ab<�WZ�8!�.�A�@5 �}#�-���;�$%j"a�%BHx�/f�ƛ~�B�0�j`��e_�49 ��\I��y:����oř��tx���ƺ
��/���7,�AY�*��3?�ږ�ց��]��~Yt�՜�;[z�ȑ�!k9o���Ԛ	92�G�@�w�MwL�"�+�� �.Mhy�3����갸F�ϳ��u��KG�iSH�Z��o_AS��]�����|Y?4��%n�wA/�m3�=tbכ������.r����� �S.���z�kԮ������Ir�N�a��4�8�i�#/#c�S ����bs�Tu�]�3ش0��{K���Z��/�b�!�f�TRfs�����Mf�g%=F/cBҏ?>rɲ����=�2=n�W��*M��T��K�gQD|�}�O����#Vʆd�
ӝ�G�8�!�8�ʵ��Ҽ)*�ҽ�T�tXUX�8._�8⫹�8Ao�&!K�6Od�;�ߘi&%;���� &�y+���]4�ڢ��)�$���[8�!�B�\P�)�l�k��~%�ߞzB�;�3@Ju:ܔ�r�c��ai[y5D2��^@Y/�����C^�xg(��:s>�MC�d�{����R���l�@|X��/�s(�ؗ��޷����}.{ܐ|�69Q��C�h�c}���m5d���D�oZkf�!�������mbA�k;|8J��КM���)h�%�I�P�턏>���Q�Q�����4�l�ܑq��	��G��۶���;iRC��^�QA����zD��}GE9}���P����{D�F�`¥��eB{����a!4��|+��7�,r�Gf��|����!C�� ]���-�k���}�,��lb�?� ���r+K��D�F���%�_a.�oo-���em��O�0�7������T�K
^9���⚰��@�I�Ot9A�;����LL��fٱ�����巖�+*�u����d��l�u��[&��T8Z��&𮴛���N�u��Ut�M/9u�Ph��v	-�N "���z��E,��݊��Ո4��h�
U �eyd�'e{�!��8�3�����*��jYYTY/�0������A�+u>
AMՄ��+4Irm�o�����Ar�1Z��N$�����(@�]�˧gi/D��؝c��j�^�����]�=ik�9��p]������[�ln�-~@(����5 ��UJw�􄩮B�ڋ��:����]�2*�@����Oナcb� �'�Y����Y9b̡���7f:�T`;[����v)������x�к��$1�S#v<�!n��<�4�l���2��4�ޜ!�Z�Q"㙲��6=�3��n��蔠};^��~��g�H�-���t��\E�hUmA
L�o��g[.ݫ��S�]�/�Rl|J_V=!\��`L�6�=���܁���ƤJ���986Y�H,����:�����X:��\6h��Ao�k��z2w�tyS��O]�E^KۺP��G{����8$|.WΤ���4�[���^$���b�wD|���;�����q�T_bk������d�P@T�|5�a����(r%p�����$�T?�|G�m����t��BL�C{pwЩI�!;1��Qr���"��1�D�+ʂ	��+�\��{��a�H'���Cg�e.�������{�33����t�*��$&&��Y������3�"C�s=z�w�H��_o����يwo��g�N��Wh�~g�Bƺ�9����0&��7E�B�A�%岍�ս��:������G���7Bw?H#紛� ��B��Q. fo�f�8�Y��P�F��΅��>�Y�:���i��2�s�����vO�a�b�Ņr�lfs!H��=T�)��>�5�S��+P|C�6:=�J,���F}u=FIYC�_[x�$�7P���o�E�o���m�R~\U��佁�g�u{
���."��_�/"ɮ}��M����+e��3�����Ô�o��3�&��=�5%��E�j���<��w���jq�t?icf�o�vmԶ������MA�LX&�� �[�(���oȋ�
ʩ%�����ņd�:��:x� ��?s���*([�&�4���5�x/��豺�O6���}렭��/nAql��v���� �y�}����`&�i1~@=�$o�d8CBV���v۱5*84H��Jj+��eM酯)���"�ap�-6
�n���83�	��rb[R�A�C<0Pa����*U)�r:��2����g�S��K9��U<�G^e����c}��<��*�O��N@�O?�\ĐyC�]	[XFz�RD�N�h��ٲ����p�T^�.�A6��A�����_�B���a�t���ѓZ����r�f0��Rf�-v|�X��9ݓV9���ֱc�N�f0:/T��B	X�$�T�B��9[�im=y|�e��6� �����a5KC�H�'�5%�l��F?-�l���C" �ө�l��,��+8B�,�f݊AI7����]��U�0#-U��0��5��^�.�Av�T� L�m}��3�̆��Ւ��e�ꖍ�1ܣwi~��C��%�wvq�a���Ϭ�Ȥٸ����.U�0����<ΚB_��ª�t��"�Y'�F���1'�)�˪ \�,z[Cg��u�` �2.�e��	��D��;9W4N�qq1�siɚ��RB��''��B�*&T.�\h * �}p��>�o����^���t�z�(��:�Hy��UJQ�Oh�����RĽ�O�yUв���3s��Hژ*��2	�ϺJ���<�&h��Oר�V>���J����rԫ)]V����=}W��_��Ifo��93�l���ߘ��oK�S���)}��-M� ���B�0l�M����Ċ���V���}�͟������:5I�2�-*h��V=ۭҫ;����BWq�,�!%#�KC����g<l[5}���{�k4�Y泂�����/���b�t+�5V])o�!�����D��^}�i�˸�TW��t����ѭ�*݀IF��!j�