��/  �}k�nϹ��)'d���V�Cx� Z+�g,��|7�mE���NBr���*��s=�M��A��4���?�
�fp���&�9FĀ�4��[Wވ4+��(��W1_�������6��9�O�CV��"S��� ����������R�Z���JI�O�����'��E鰪�!^�0d��o߹���ɯyw:=G�`�9�PyCE��8%X�7	]�*����pogU��(~X� ��Vrv����P�Uh:l���V�	�$���p�2��_1y�ȯ�u� 4�D�M��hݿDI� 6�pn�l�!`' ��-1�=<H_6�n�������@� 0̦�H>"A��5�%Z`<�\%�v��>�cy6�f����^�)	��}#J]�/Ev�rgQ���Ըl�S�%�陣$�#}@��l�7���w}oB3���5T�M��ĳ�]��U��ɶ+��t�r|����az-����J�f���SWǦهK�y=|6Y���ڌ4[�^2mtP@-g�<�.����E�To�ٷ��ts"����9 	<��oؕ����	����f����ܫ����*_9��!�7�R/l�ׅDۿ�o��Yx��LR
�ti�t�.��S,,h�f�q�����	{P�ȸ�\�/���x����h�jT5��G�X�"iSCB�R��Q#���J��FI�Z�?�{�F"�H���^pQ}Q�ب������4Y=
D�S�"������@ְ��>+@t�/�qݺtk.+�x�R�.�PJQa��"��	��Q6��/,�����'%=,8S;"�,��]���^���nU�%�.X�\)p�n��bx�H�¹A���8��܈"0~�V�SU�T�_�eܷ��(��8�������:5���-����1Y�$�b��)9�oQ���	Qg6a�i��B�bZ�i9ǚ�^4(p��9�� �'��|Y��­T�wJXЪꢡ�������x�խz�ԧ����w82L?���֦Z��-8{/L�3�5
�,`pI�j	���`��o�c6�5�g�r�^�Cr��>o�m�u��T�#���uB���x���rF�8%`r�o��0�1�0����.]F������)~���&��i�O�p=�p�䕣��G�Ң�G�r�\s��J�e����y�~3,�pr� iُ��"P�
�R�;!��r�Y:��G�-�$w�1
	.�c�Q��F���}�����lk�����s�I�x魦}��4{�Rן�%�{����c�G�Ѯ������W�s���pS�.�ͫ���Tr{v��z'"��X.�s}:��l��k-�z3 ��,�ٴ��ܧǳ �J�3��}��9fI�_<�n�CB4�h��~��Ν���N|��"2��M�ub�ܝyW�<����( ͬ�
G�ϣІ�$��3����Ь�;���ҡH��C���(%���{���=y�@�:��ϩ-��z�|�d������sո`.����L�^>Ǯ�hU��*�r�6~�[ �vo3�C1r+4���M��Fˍ�d��Cv�����ԇ���TB�K��������ۉ&��:.^�.-��aݔ��|k|�����9�w�-^��6�LT*1UbCg�F��}��Y���sS�LcK7���I�8����iB\�\�ۚ3��OdpU7��23!�������2�l���i@� h�VO��8��L]��(��7�W���D�D?׸�g���Ɏ�=���&Y�N��v?E�o�S����R�LA��
�T�~0�=��t���>��S$�@�M�����Z@m.gi��8��[�;xɪmަ�Q(䑔�)V�����Ʌ����[8�w�<��z�Q�_��:��]1��D}{
��ժ��v��/G+���$�w�Ӗ��>!BiG�̼C⚪[�ߦ$��Y*f�̿��98_��=^`��E��d���{9'���2��w;��PI�$�0�\���\�S�� M��p'�-k�&9�O���x�>�1;���N�����N��#|l"�u�o��=o6�Ϩ�a=J�R[W1彳Ro��l��B<�$� �Gq'�L6p!y	���:Eڽ�B��[��NG�F[�����V��Vj�v(�gc+u����a� 2H_���R� �_������K���G%a�L�����Y0��������=J�D3~�k6�����Ãΰ��4C��Q�y�.%p6ޗ��af��Q��M��.��&J���r���퟈̃���j���u�:V����N[�w��_�q�J`r������m�P�}Π�l��	cNg��uT�g�[Ma"�Х����T�rw3ᐠ���p�߄,g! �a�9�u�U�)��>�̲��$��7�J�����ld�}��N=M��ؙ�nF��=\��F{Q�$�2Z�G|vΓSؓ�0��F