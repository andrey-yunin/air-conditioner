��/  #y��W��K�\��H5���H�=�������N�47Z�Tn���렙oq ����hgg%D�MБ��y;=.��i-�CIEO!W�:��m��M�&�{����e;#��a����LY�Z׷��qƲu.���� ?lf��.?�W�<�"�t�A*���u�簪�!^�0d��o߹���ɯyw:=G�`�9�PyCE��8%X�7	]�*����pogU��(~X� ��Vrv����P�Uh:l���V�	�$���p�2��_1y�ȯ�u� 4�D�M��hݿDI� 6�pn�l�!`' ��-1�=<H_6�n�����ã��~�������T�\ҭ�
ry[�o#�D�4WO��U�}�o�P�T�cbT��d��\ר	�km����ܷ_� �U���uM۫�@�`�? �oPmԖI%�(��؋T���|��#�۫�bΪ�h9��T�Qa�n�I�ȼD�xT*�>��+�v�X��P�[��,�5"2�����8��-��j�bB�������D�kE�5�ޕMF-%#�z��/y�������N�C6�ig]*�vl���3%��Q�H��('XѤ�V,VL������7j2^V�w�R�v6�(�\D�WiKwo�����shQu4�@u.���v��ߒ����3��@,��9�f��U�j���V�`�>#��A��"�I���P�u�5i-upX�3�)B�1�f�U<��@�L�H���y�]������-Q����2?��Z�	#�{кA� �b8���d��~������KQ�n��c%�v�f�}x(�3٭���nE̈́�'c��n�0T�ģv	k�o�_CԔ.�@�Ԇ	V;�)��N�P`�]�ŧ�٩�We�U�b��$���r��H���"��B8��Yj��ڙ4y��p��2A?���0��u�+�ʡt����x�r6;&V�*�5��P�s��lj0��7τ[��W��p�.
@�4Hp�1��h�,
]����Ѭ�),.�G����m�,�)N���M&�5��< ���_ӯ���1�m9�:�'�8�#���h�4s�Z&�ΫC�V���p^�F|������c�^�b��^�w�cW��Sھwd�yBN���1})G]_z+w�n8p���u:�ܿ����%SJ(�����ʮ#��U�l5uM�K&�Ҙ�{P��'�]�n�7��
s"n��n��=�#<H�	mV>�*�V~�C���. ]�b�N���
7��Ì�m2��xPQ�3�)�V��JNI�Nfz�+:ci�b���^�e��R��:0�q�)Bw�D@v��>Dx�~�9Ȧ�;\�
�6*�%��U�h��j�=�=	va�������;g# �+�y�p0?�.�{ZFH���1��w��EOJ�fu=��h�̺�g�T�_]#zYi=Ჭ)/B���4݋�~��a�G�i{N�:�G�v�����lg'�%��3/���f)"�j㽉�@�u��*^h,c���fk��/���jDw��:ȣ����.��N
���l1�����2No+MwS�������8����9�n�+��2D:�,��/*�1i݁���Km���V#�`�	`pG6�O~iĈ7���.�2�t6���3��{9�;�a��b�mRƤ�>�c���Pɗ�z&�p?)U����ߴ$.�1�e�n�bʩjC�Ī1��ae���J<�6c������zF�$X��{/��$�ٍTk3g��&
�mC��s1F|ɥ�/�Md�{�]�Y�P���h�<�T�4c�OG���g��zL���x?TVD�eq=r��n3X�o޺}Т��J!e���Z^�^�Nj�!7�%CR_xzw�m�^�� ����f&��G�#K�H��Ă�5eDC;���ݻ?���2��i�Q�Y.f�����B@(����
�@�����r8߭o�j_�C��U��xE��˂��n=��Jl9�x�� �w/����΂o�_��A&3���h/�ʭ��d�-l�%bԬ.��O?�l;ﰶmj��a����k�@�;�_lx�U��>�/�.$1ybt����t�8Dl��dTS� -�9^��,Ӈc�ЈâzUw�T��W������m�n�R�LҶ�%�%ϐ���_��D6�V>�9򳬾�	e28!�Ԧ����������ůU�������?���"���V0�����* ρLx��$G\٬�j�j{E�K��ꢞ;	�=�� �j̶�xp�7�G��GC�?��x5jbC���em�������׌�����ukJu�;���+E1�������Yf����"K:~��H$0�\s�WH�R�-Ο=B���Cn�~ $6ExU�����M�F1j[�nṘ�/XCO4�'/�NO,�hxB�dqX2b��;E��⚫li�bW�����1$C�ԕ�����V�;T�Kp�����x���0�<3b���	 �٫&��!�C[i���};�qa`в�&w=����6Z�K^;��o���k��KD����oY�A�<��E���YRm�HQ򜳅����z�����"6���@-����m��K�� ��O���~!Ў��ꪟ9�_JD1M�/(��?ܹ�ș@J[@[4�O�D���A=0B���8-��zoL�
�� ������5I�Q��g�"F��jh�� �FIbU���8I�tZ�Xz�Z+�_�xw��r���ZP��(���"�	��e_���zLz�8�ڋ��,��_�E����;��Py@��E��&���	�?4z�-3O�h t��R�F�d�p1�z�`#Rau�'��.NΑdG��{v�H��A;�X����I��/pi:�d_�>&���GEy�T�Q|Ik1r��J~ϗ����Et�1�l2z���⛲I#��jb�Y��;��'�h�J� A�ۣ����^2��G�p&"��|Gـ`��Λ�z��X#;yr�JX��r��d�t���uv�*z�V����|85�r+��J�I�,0CU�B�Kb�俊���UDN'��\A�`���P�����[_��F �w�`k08^��dIȆ���?��>����ՃF�E`U�x]t�B��^�\�������j��8$e3IJ�v�^y�A�C�CXp[v�]����2�xOJsBCnr�dl_�\�:Vf���=��TXN���(��	�S�>����՝���K��-(���b�p�.d���z	-[v�@��9?��Fe8���ҝ��T��8Y�=���AN���P�~/(�n�W��.�
��BǱ�s��g1Z���	�rٙ'8�U9O����R���Ѐ�ߕ;"�� ���*c��G�[~�g'���#$V��JR��i����Ε��a��w�]��XP�g�ZF�ih�bʂ�/tm�]�6���K�dT��s���6�E�l|�e#n#�YW������.7�`���-;��C��^O���N�Ma��d��q���8���^��ѯ m_K��Z9�.s���7��=#fĒڨ ��h�t[$��E9�Л��L��]�/��^ 4�[�y�*�e�o��X`Ԝ�H����bAA�YK�7�۷��#²T`h�aH��J�e����6�Ȕ*�*g�p�{�H��t�6�u��T��K&?����^�d��!h:y��f&q�F k+W�ƨi��$���1��E~��4,@��`�=�"�����;���cOx�$f���1+؟:qT5���Sɣ	������^Vk��,�j�"k�����bZ�7�K�z�U`~��+�������\�o�P�(=D���Q�c܂Ỉ��.E���/uf{f[ܺK����(��m,��K8{d=k�Ixt���xћ���t�n	�!`�M�n�C:
[��b]���L���B ��U #d�����r��bcĠ��xѭY��T�!�Nu�&�^���r?�\���*����FX+]%snp����c�V��B'�Mmi�Z��לP�1:(a�3��D�%����H$�����^�N��U���0�t=��G"2�䐘�\TQU_�q
f$b.H[�RȘ�������V�����Ļ	��6a�)u��+�=O��8����E���:!�+���;��v~�;͏^�{v�`�B�s��?�Fj5�f�v|��,�
���p�ٛ�ɐ>)i�0O�<��v�ڎ����1���c$5�����O���wo+��$2#HK~�ʻ��&ǏG%���(4�K�[RD��x����Q,"-?H}�@*�]>��T<��܀~�f4��sd@V1�19,r���ꫲy���E�/�rBo�N.��5���
��/k1Q�b�j&�w��
��4v�	�(Ƚñ�$���E"��(#�qR_������2 �6dn��I���o.g�<D����Ԁ�+ll������b����	J��sg���z7_kQ�tH�����n�9��'ML$��l<�Q���ǟ�T�z�@�L��l�nW��F�0�-(s���,�2������?�9�;p[4O|��tu{�]��$͊��d��܃PR6"{���.Y`P��}W���@cM�ڶZ�|vV[� 'gO-%�h"�޵�9�T}0b�7����3Ar|)�S6��l�V�n~_6%'���1�"?Q/����$�['
��R���#�ƌs�^ x8�#�U:��u�yz-ԟ��D������_.6́�$������
l��Ҭ��Z`��0�4��B��>r�ֶl����M
�����u��n�/���t�.�hwq�&���:-��ERA�{~�.zFmqU�K}׼/*���|���Q�ZȲ��!=n�'l�	��Ф�%�����y���c�:bF�f�d�W�hcA�g1C����O8ߤ���4	�\�d�KU��9j#���>���V4�Y��� ��ʠ���	U�����[��,n�^ĉ��f6ˈ����܈ɝ=\븙<�s���gK�LJ|מI	��dr����^���,B"�ø�}�юr�1%�Bw�4���l��w��,�WA�x>�7>ک�*��i�]�7GC}v��N}�,�D����w�1��j�%�sQKP�1ڮW��h�9�+Ewt��AH�,� ��-��X���ւ�ǅ-I�i���{�Q�F�+����K�5�Jn���/L�'J���TݩO�.��vL�s�@�̌�zEv��$���?�2K?�G[>:����q�$1�t�dG��͜oyB�VL=���C��y��<�d�5v��.O�\(�6Y}����G%��tF��\~��EQ��M��d�Wa�x�K�ј4�S����8b��j�Lc�8�蘷�x�\��8e���z�ߪD
Z?F���S！F��-6��zo�3d�c%�J�-�@��������jUTԂ��`�rQ�e�X��~#�U��=�%d��Ȇ����=��oҤ�頉���e]�`B�z;!U�	�d�n��*qW[�_hT#��sC��Yp7�t֤*?���^4US,��>2�I1AG��/��v�v=.z/�ݞ�w���C�O	��W��&����ܖ��?n	}�հ�������|.U6O���Fb&�R=}]P�$%�}�}�
qq��H/��X���&p� �zy+˯�����E-��n&Z�O�b �_�o�՟W��!��D�W�u����}�Y�H��a������q�m�����q��+���?l�f�y�X���55f���]`��Bf�2˵�Mk�����d�_sÉ=���IxN6{�8U�ȩY)��w|Q_��������O-�r�A�VWO{������~����]ېr٪{o�4��zx*��^*XяW�s��~���8[�/��Q��8y�X��.��;����؁��w����;��G��W��#�G���9����7��;<�T>���R���5�����a"g����7ݩ̗*m�B}dyo�p�Tɾ��]9��G����M���{��ڽ�N�C�SbnރF��î�M�>a�h�En.��99;��1K%<���=�k)��̍M`NڎsR�IwA��lR/��M�U{OS3��J-o�ϒ��KTK9P=T<��TO��ĉe}Y�
�&:-��ķ|����8l����TwtV��5��H('��x\'��!tF]�и�eŠO�<C@��A:��K��dH[Q(�-^�>����}�Z;�'7�X��n��iH�J�Q�d�ɐՔ>�<nVk{�7vq������E|�ZA�i�Y����c�;�$oВ���RBꁎ�h�2'��6b2���擈&z���T��q���6���������"ש���q79vi�ѩ\OrTi�X8�F�$,(���.K?�h�46Is�-!,F1w8qF!�X��v P��~��RZ	�@�Qeί��Z��7�s�u���H ��-�� �H�X%9صFW�A2"y�������1�q����I���� Q��`��6���,�b�\��Aw�N&͵��Kf�?
I$EA�Kg
z����$񸫕��
�֘X왶O�eW�"P��]�^_~^�:��.�[�� ������G�N� ��I�yɣ>O�[�Oz9X��(�
o,?���zN�Cu�0� M��� ���y,A	n�hpR	L��E(G�C�}=�w~H�)���J�=,�D�_#)� ��f�,��o�F��u8Mg@�(����9��
mB�c�����5�7v�bc�~6�e��6�CD�=��_��pǬ?3d6�ʕ��yfh�R�MZ���`J��͚@��*0@�f��Ÿ�!��)���[�m~hj�u-����'�f�S�F��΍f��t��:n���x�����`�w):����P[Ż.��W7Y9�ڔ�Dv�L�̩�kO�l�.xeEG�`���z��zȲ@ �Lj�����4�Ê����\;u���p��^��O�j*�V��V@	]A
��c�#�����V%aV��&*u��hKf9r������0�I!��Du��%wo��GS�Pv�k�R��y{	�L�̥s�e-��۾} ������O�'�n�\/f�d}��	�*�^TO���j�b�oe/�9R��s
��E`��V�i)�Vh<�2Iv���ِx���O@�F˝BjܦT�)��6pm<'G�ɚ����q����g�]Ή��./�Z��<b=7M��t�8<�m�""iW�@sM��l�� ��0��j�U�v�M��	%��{ҝW+� �H��h�T8��_0�j�j��Q�,s{/W<5	��U��>$�_Lq���%�SxyI\�_B�a�u�"'0��2��D�����Z^�3�3�~��m������9'd���ނ���w�!���xmW�%��t��J��#���J�����1/Q�t:�<�]�J�.~��m�؞y�i,W�.�k*M��e��]A�m��>���?d����6� ���a=oZ�K'1�Ͽ������K�=����C�IǡUV7����L'c�V L���LQ����eju�C�(j��0�P��{��s[-������O��#l�d��ԆG�o!��o��1�K7gu���L��<%�ake�k�B��� c<k#3C�m6�g],A"��G.
�C}���0��G~�r���Rg�K< \g��+b.�q8��2�u�x��-ϐ��Z�̒��h�x�7�4\ӍMM����*Mݪ���pR)�Ǌ�\�wP±���s
�ک�!d?��f�^��.�6�g�X��]��sI|k\�r�~�|"F�= �Ŋ�wy�����f�ő-��ao��+EFT/�0��`���z��J���IO��[Mn�y+�@Be�� \q�7؞l��3���j�¿>�j������&D�uܖ�;���5!��Ɉ'�bɐ�����n��n�d�b�k��-b6����8'��H��)��b� %��.��sf~�QǬǸ��{���ztX��ҋ���K��Q�u��2��.<g�mNv����n�`�5I��q��� d`s�B����%
�� �b�P�pPE�2�+�������8�b���C�>��I���9��,(y?`ӈO����G ���_>��P YNױ��k}�J�
��,���7���?�4�i��j���֤�Gn9y�33�;^��S��K�W�WNv���f��Z{X�,&��p_���֑5ay��&h��|5_|���Z	,�xS&fd��w�33	��m19^"��J�N�@P
lt�)ɨ���6�s�n�/��0���O�����m���8k��A�fr�m��؂�s��,Gk@�;1x�� *�#\� ��[~��ۧ�6,���k��θ�S���&5�e���0q13������󙙪�&���֚������ �áa��~���SX֥ձ���r�ce̔��!p_�rM��Q�jtE(7����!�C�[z3v�I�M�b�����2 %�'�~��"
w��;�.��_�/�bp�Z��WPjh���a�@����[�ӵ%�1>4u��P}z  p��YQ�W�T�Ԏ� $��	_?��ww�O$3߭7�b῟W �M��U8�r�``�e�Gwu����0H3��E}�ش|���:U���]��n�qSآ�/A(J��OWY��Ԕ�.�&~�G�R��_g�/5��F�M�3{���L�>0I0����q�&싋�8�|����r�L�r�8 z����v)�T����M'KS6�>>���	|HW��� ���7�ۉ�7�XN�Q��W��${�Ui��wQ>(���'lf$kP�0�qmց�o_��c>�)�|9�2����݅�a:��4N��`Ҭӓ��\�����Rȍ�D��=M��Nh<�Ð��y�_����%Q�Γ'��$[��M-z����6��)�*�U n�x!��F�Οd10߄��n˾cնh�3�1�pA���~x<�H��=T�j�ؤk��c,�%�T�TiY�b�"�S�4�D��i_�d�IZ;�,��}PN��ݨF��DL!��j�<tԐ�$�i=i ]�e�b��m��LO��ȸ��b� ��e� ��ğ�t���8�A\�Q�zW��%����E�Lh�{
<����Ê�F~�h���[�X�U���{ۛ��YM�b늟���pf��TV�s$���ϩ�H��U�_�n�v1�^���&�]�,|���UwX7�Np�L�<u-dP���zl�tr:ŕ�,YO?��9��ځ��:�4�a���1R�7y)������X%Fi��&���g	K����N0�)E<����!����54N]�}�B�F�o�m<]�7|7��
W��?�`O�I�0/!��y�C��q\���q���Mޠx�w(ƹ�r���}/�'[;:�M{��
|���ʹ��"�.��V�L,ۑF�%�X���,v}k!�`�p� ����!l�r�( �?����f@Z��N��x[����9�ý��mD�~E_=Ӛ�I�)�Z+m�P]�fi�pw�͏T�^��V�v�5��X����Egڣ�MpC�*3�!�9�P�چzE�q2p��iΉ���x|����2=�;7�6T_f��ί�Ã�Y�{:2�[� �������*��V����uzI�z�W�&A��	������{,$R؋�J"�=�[\�߯F'E��/�Ư	���VVH�s�1��^w��	��dJ�s��ɟ���\"c�����1»��a����j�"G&��@U&w���-Zk���6-�AS3`�	�ro2��H|�S���E1|�t��5[#�$��/t)ׁ4�p��0��� �ߐM|�OGR)*���ć�G��~]�ʳ7��;�����{��_C2�˴R,��YB菱H%�.����W��Lt�'x�@�c�R_���`��o)Zs��ؐ��R����S��Pt��76�*��� obOեf���;'�I����`��v�~w,���V����>���}�S���Ư眡/�yj"S~�����!m�?~���Z�n�g7�|4���<� y� _�E�2+@c܋��T>��6#�Ia��O�jj��N��?��p����D/W+�1v��Z1]I�v���A]�6f���T&�^1��em)����_��°�hԈ�1��/ّ�����z6����LC�*)X\ؗP�<h��Y/!k%��SޭMD���&.�r}���E���Y�[��'�xbB67-@���hb,�*�kؑ,���ۅ����T�@�* ���0ʥ�!�J}Ig�L�m�ht��=�ptP9��n�ޮ,3��G�~9-ñ��7̈́�w�e�/q���iyA���j-)-Oт��JZ����w6�I�'�4�E�� �p�Y7�v�Ε���(���$�Za��y��#�FDs7��p�Zt9�����'<���O��~��I�'���B�>X�WG(Ӏj�{!��)�i�C���>��~��������U���o<�Vx�֏�F���kd@��E�AdDc��ߗ{4O+�ȧy-�.S�'��9 M%�6Bx������a������p�\���l22j�:��G�5&r�m0w2�i�}�����}�TZ�N�dz/�C0���y�g��'�/+��|q�+�2p�ǀ1�s sY�#�-|�Y��m��"M��ƄrWq�?I �\����}g���b���(�쀎��Lhj�9߹*+�d��,������~�?���g��ӑ�[�=-egC�ڟ0>|[��d�3��Z�:e���1�{��G}S��P!�Tڬ5^遽�Z�ׅmQt;2@��W`�1낇��~��l��QğO��އ�BI�M~N����}�Xr�P�tl7s����H��Ycz�����"A"�>F�g�?��2
���0����n�]۫$,o����j��qF���HV�O��}�~gS����-�7���~�3�>��h�خJ,��&J3n�2��D�c��f���_|L��8�݋("�x�Ǩ�o�.��d�t�ɩ�lF���]�t����R�M��M�`��Y)����F@��;��U02?A �x_���<�:�iA�xL�1@H�zp�D�z鯤�+�>����Y�$䄹�O��v�ѡvO�y���Mdq&k��>r���2��,j_v^����)ˍ$�0*�	6�ম�O�'R;O�:,���X�	���E�eGB��%n+���X1�Y-AI�����ʎTT�%u�0�������`a/�/�SRq�_A0@�::؊�l0;S1	cƸ����s�����ٻ�̞qsծ�����
��(ˁ�Y�Bb��d��v� g��H�p�&e�q73��C�G�w83�e��f?��]h]=7��Nv�vφ��b#���AXlF���������WLt!w�!0(��h���9톤�K���i�i��;����W�erʊc��·�n�\)�>ɧ���.M�����n���7�߼R%��R)l�w1���]J�~@�I�_a��dP�ں���CYO�d衔'[����ٙ��;]^j�ۏ��o�_\JۙK��h�N\�����~{P���:�-�\3�Ar]�X�²r�F���iqd��4���X��u
��[)^�*>�c�s�hҢ�i��SUO@!V"�Q�M����U�)��l����ڳ�n���V�q��J�!B]�J��Ӹ�Iu^.9���m��u++^���~����I�����{8>2@c��I�o�YJ ��MM��҄�d��˪�,�ߙU�C��Fex:j�B>J�~HvÅ�d������&��c.V �0���
�:I?w���W��/�E�o��Xu-��i��r�0�S*�B��,b\�O�+�+��%C�A�ZDa��e�u��X�9����B[�,)�����oH�����(���!�HOuϐ%�c��Y�ԴTV������V� �>�6d�qu�|�P�r���#Y��V0z�� д�!q�"���cd�#R�����h?�^�����3�9�>��}�ג��]��l:�&�8s���Sn8C�"
n4�
Ѷg!��"[�+����I��O��qpu��Ҥ(��Q�mTzk5�ly=\F�����ՋP�.�b�+��	��gy�)p/A��x�giW�(n��� �j�M.C���k:5�)�m���n;я+�ma���/�x�d��3�F�<�/�,����:G"�q������!��0���Ȁ� n���^T�8;�Qt��u���xiBʂ6�w�d�ҋ,�Ӣ7�wz���"�-8��,����:.���
�X�Ә$>����a�/�rޕ#��̆�W�����Ha$U'����$��o���"��g8��J�v;§ջ�k~���vm�[ir]O�K&�����m7v/��>,>��� O�Ĉ��������U\V���vȹ��Qn�^���-q0����=��q4I�ɠ\�`h��������E���.�+��_��7\��$��@u�&���|� ��&��%��bO�m�s�irnA8��6��ߨ�nmvQ' [�i�?���]��;��᧡LM�8<�Jĕ�V����� �:�o
-��B^�I�2�����)���B(���kI�����^E�=Ъ��q��07A�4�\z�
�'��B+H9�g?۽2��׀�u��\ֺ�j�;+J\I4R�¥K<�H�u�����{@,Ji���2��� Ve�h���p���%;��J�˽ep7����y�e.�3�U��	(�"t��[���d/�?kG
I���	(��^�Ô/�"��pa�>�2�H��Q��Iī�(c�S�2U�b��L�c����&�3I��h�5x�  R���q�F�=�����J>h�n��G�m��܏
G3+u���uZ�C��F#��_�Gv6���\z�C����]�j��z���OZ���Nc��_QMr����Sb���TaR�'WҟRmd���D�� _�O����y�`建t�׫^k�b���?2�-9@��k�Mn:�̒
^~�;�Jf�|d�=����qﬄzj�����H"nZ���YϭyIK0eݰ��~�*����I�ϪBt���'�P�mA|)0�ws������8d�Ba�����fW�	JsH�K@�r�]���ݣ��z�7G$9�)�A�5v5�T�9�ʒ���C�ɧ�x�C�_���s{�'ː��R��+9݃�˵9�+�e����ݵ	m�F���-DxH�͢��d��BPM\n@�DwE+9��������hԗoW%�q�u����B��\�7݃rq�x"�N�l�L	Z����S��fQЦ�����9aZ��i��#*�m˃x�`sˍ���A��
bH��e	����-F�^D1K���T�t�*�����lץ�����SH'&�ڜv���۸�(�pm���zA�mrm����c�wl�@"�Ӹ��~PY�m4��h�8$�*:������+��z)���Pe8�p��詘T��O�݋d��%nZ�� 
�K�l��t����m�.�&�74�o����a�ϊ-�����jm8�k������������AU���=0W� �������J0۳o�<�
��Ю䛼��i f����'�2�������%�Lc�Gc5�����2 �Л��:2j7�]9K%��
~Rg��}"u���o��Uˡ��3�_^׸g1�"��ǅ>�p����IlmK�	&���� ��q�3��ڨ&�SF�aU+���hS�'e�
�����?�"�����9���NK�$
���@'��ȼ�},�{�{_�ˊ���� ��		��z=��c��I����m��#�Бb���"k�[�`Q��UY��c@̝�2�7	SP6s��;���e���;��������$r�P��&�(O�о�V/&p^�,�I<r�`U��d\!��XF�@%}�'�>=�q�R�EPL������E�m��!3@�sɑ^>��B:h`��W�ó#^��|�ț2՟4��]�Շ�[��D��C��fY�IH�8�avO�2�0�S�Zf�O5����1��*�2����iP����.��^�І����G~5�tvA!��6�*�ܥ�Ic(������%_C��tr������q�摕'��da��vA��Hg�����pPћ,�����Ժ����^��CJ��E�Q>Wf	�W�h(���3��X���;n�ҫ�K:=<V&\3��t���7�^�b5�����R�~G⯺%��`�/��Pk+?���k��M��^w3�#+��)�|�Ԥğ�M�a�?�#roV�Ly�2��(��7)NB��BQ+j
��+!
�~)�x5d���ƞ��k~$��ZL9�z?���0x���TN���ڌ"4Ʉ���'+(F�KK�>Ċ�c���ka�/����_?��P����{�gj5w��i�� ���
p:8�mQ�E��B��7�<Ғ�j���9|���^6@.W��~�~���O��{��D���y{k�c��{B�^�Wc�2��i^0R�b�{�����̝����,��9�K�_.g�É�1ԋ����'~�Ǻ�҉:�G.�#b�B�t�t:�!�yZ��O�.��.�(�ͦIq�qM]�Kr�kq�3��r���S��)�o��֓Կ�Z�<
�� s�t(4]�4���`������[w�8�O��UxB�9�'��eqI2��sVO�.gQmp���o���J@�Rv�w`�ة�i"C��\�|�'jB���sS�I�n"�ƥB����;ir,6{Th��MDJ�_�^�T���_J��;�a�� ��%�a��Of(��	�>j���θT���t�ײ@XR��D/��!��^,���m��הM��֞:�-�Ѿf���.��]��� C�� r��ퟌA�:�n_����k��e?�7��J��G-�g�~:��QtTI���n��8����ՎHU����0�t������B�L�f&e��I��Z-i��Kx؊L];~L3��t����+����9O��@�laeHi,6��W;<#͟i�}��xJ�C����񒿛�7P���N�H�.cxK ��33CHV�<1��"keJzb԰:R����N`^�9r�ɾRQ����E�v%h`��Z�0O��^[Y4(���Tf\�Z����'.	o�HR�S�1�y{sWCR���dv�ᚪ}��P�6����I���t)F��4Ӟu�Ft0�9��r�M���_���ܬbv�Sϡ:��~Љ�T�
��9YR���3�T��
meI�q��u�D���3�G:��~�tC���|:��§*a���󞹹L:Hxz	\ԽA�!#o�ϛ�<0�I�G,�Ҟr�#���z=!��:�K�LgSC{����Bi�F�����/,�� �g��=��y�> ~��E֤E���z����9��7�x�y�^'�C�zu�~�-Ru��7X�pZ >˰QG�����6��P6�j�9�Y~��Ӱ<�o�!����_Ȉ!�������M6���m�_�&�[����rTw�Ƀ�~�(D�-7ac۝V��ʺ~3�J�f�n^[�+�`$'��sS�9!V��֨r���Pa}�-�Ƒ7���v؍׺U���o�³~��7��l����n�y��f9���l�#o2�L9�K�H��ݮR�'r��r�����T���1���(���.o)���Ga���I��D�U��(�\f���m��6!Ř��k��v�7�UY);�[A����*��� CXpfm�>�c��"��� �0-ݽ����T�KH�x����7�MGE`���w�<L?z1}��u��3��<fRk���E��l������G��R�T!X�f8F�a���G&��V�<�C��g��Y�(���8�nF�I���6OǱE�Z���tY�]�`L^2�Pk�m��w�11��&a���������v;����2 �=�Q��#���^r=���3M���;���X�ܓ����� 
�ɥ��H6�7�]�̄������R:�$�����x fO"Y6a����H��6�^ĭ�ܠg���5�H���,g�%�T!ڊQiz7�����)����=��	^��)��� �V��^�AJ���l���ڽ� �_n"��gz|s9<�^\`�.W���%��j܊R�ڟ�7A̽�:���}V�ǳ[� XY|.��i���?�n�0^�p��u���N)����]�Q���\���=��t�ߥ=��[�f�5�>!��;�A%Q�W0�:-Mވ{�K:�!�Z]hF�_�Σ����K�3T��4l�l(�o��^k�?g<��8��T��hB_I�T:&�NQ�)W+���]��h�8j�2�o��,*����4&*Ţ�S�"'�UQs��I�ܔ��V�a$����S�����J��Ud=`���qG��t�h�9ϟߕ��/h�o�ZVt]NʸW�.�(��?]�ƀ�!�+��d������&@����ˬ 3%�