��/  G�������z������F��� m��7ў1�F)�'����p/@�����Q���F��p݆�:�B�m̏�sf���	=.7��$nٞ(3��l4�ߛJ��E��<_}<bW�N�!xoL0��E7r�DPȟ�b��A�ŀ��R8ꪭ���!^�0d��o߹���ɯyw:=G�`�9�PyCE��8%X�7	]�*����pogU��(~X� ��Vrv����P�Uh:l���V�	�$���p�2��_1y�ȯ�u� 4�D�M��hݿDI� 6�pn�l�!`' ��-1�=<H_6�n����k�u\��FC/���"���<g�S�S��S��u��t���|�@�L��>w|����\�7�}:@����Fj���Ʌh@�۝�Q|p����j�N�d�Y
�U^��a`�R�?\����3^0��o�����y���k`��&>���
�D�����-ICD:���ғ�� >��B��$�c�Z�%1Н m����uE��g�)�I�F�d�D3sɸ I<��F�8;�����r�'rf���A���
&j\���s8����� 1�^2`��� �d���1*(�џ3�!J�#����/�ɎI!�Јi���筏�Ф�y+�	f�q�x����5�&�C7�Ls��yJ+ ` &�����b*#�m09Sj�@S�U������܈]0H���rDCSs=�My�v�C��k�㎜���P�Slwe��4}�yzì�,@S��?*�i�����aO�dH `�e�]�d1�:)Y,�8�o��^<�&:�<�tU��DV|�pu�6���2k�d�������?�d�E���$����P�ګ�kl�5Sc�n�^�/Z�	���!P�� 
�7p��S>���uXF� 9�Y6�9n�Ucߊf�C3��ϯ�UJ�x.��>}z��b��_�=�2���L:�^!k9����po���J�"����*�8E�̴�@f�1P��[�"�n�Z��B�m,��6:H�koJx!�bs(���Э�{�`_�mh}Ŷ�3�sL��a3i�N��01�d8L����b�f�Y�ŀ��r��`̇�����"�F����鍄>F���ڛ~)U�J?
�'�:��bܱ�m��l��^�{ހؒ���=j�x����I�+BE(�c�]�=?b���mʵ=�z1��jx�⋙������^n�Y�����Y�/Ѣ)�R���d�喸t�ǚsO�s������z��$H�ɓ͒i�D��a��mH�n��+��Cze��퓮���zR�Z��`!�x�{�+1JʱjF:�D_2"|mD���l�o�w����?Der6+��#w���oוp.#�̸i�Y��$9���&��S-�� ,��$̾!.���>�ڴ����4���9��埐đ��Q���p�w���(؛#5P6'&��B�ű~��oΊ�;3UN��:�:���?��ˈ���C�N�����x�SP�"dq~�,_�$,���%t�g:ɛL��J�L�2�����Ý��wZIw�@^'�Eί2?�-W�"��N��6	t�u����9	O?�|��+��3���b
D�-9������b�B�9��R4��v�;m���gm@0tCug�	�(���fJ��������(��-�X�h(�L���^ĺ��H�f��+*��˕��P��@"F'r|��I'6X{3���QI!ܥE��/S49|��R@�>��˵�zNץ�ܓ݇F�;�Sw��κOsW�ټ�۬�L$E���m0���"9Z[�L�$a���f�D��@����z��\�KM�'�� hhJL9�`�>��aQ��CɊk��C�����RGI��ޑ%۝5<n1�KBG�0JQ@�x`4�R"�ꂻFUEg�B.�ߥ؅�����(C �f�QPי����U���#o�>}5�$-����s�'MO��^)~O߄x��B�i�BH�(�O2T{ ���i$��<V���A?���Э7>��+:O��w�1_!�A�H`��m�~� �qB=HP��͓�u6�e�;AH!N4t8�p�'
��U=}nTu%��.()�.�g�/6�:Z�����@��҅*��P�_���ʰ��=�)_�lq@�����x^�C�=	N6�NI7��b;S�qx�nS!��������D:C�~�Q4�;�c,	�lZ���q��jk,��JL�3;�����f�u8��$������~��H�r�u��G?$��_��_�N�P�v���H'Z"e�=k^c�=�x��@'�WN�I4�Y%���ajw8��nj�~ѬXv��U1�&�e��qn��V[#X���0�ȷC��B�gIZ�����8�v%�)h$7�O�d[�Go�����{��&��-1w�:½M��Y{R��N y]��&.�thlNv�&�w�$��������J`���@{�
^vBϝx�Ak� ��~+*9n��%�����˜��*�i�ֻ*H߷�$�"�ǖ
1�JJ�+E�8��"yZ�	�˘9��v`��|T�*�D6��5fa�69X��TV�� �z��^ �e�/(lZ�(9qH�����"o1���D�{��~ڐ&�e�j�e)�^="�Bo~YS*b����5[���6����0�g��0W����Y��kh�#��m1[~�'�}"�ir��o�=�:y��(�t|s4��[V�u�����҈�"���)�XUS���1����L����Tk���Cm��������E8�g�,v>�<�>䉈��ҷ��A�Yh0k[�}�)�Aj^���A����7?��n �&���V��(��逡�]�X�M�d�A��vH8LZS(���l�b�߭�}�f䯩���H7�sp"g��a���*<�Ԟ�w ���]�Ř�s��eoe������+T`g�Ű���ŗ�_�J�=Q�ą�y�'G���*�]����������D4�QQ���G`��8�8@�^�)ExZ6+jw�%��2���0�au&|�u�M4���b۠?��<�(V�|���S�r��Ķ�J�|0���<��jUI��a�R���<��Z!���&7�y�f}ж����)b�ܞ�5���{0�D%�C�������x�-���4l)3� ���O��Y���ć���e���v%7��H|�s-�j�yM97�q���������O[�,����s�����h��g����6��=r_���f;�	���W&�q�X�.G/���H�|�9uBwt�:at��[���4�:�������V�Ƶma�#����R�!uo$����B/���e��<"z&A����v���tcӫO�Vu��e�tŗ�1�a�����ЂO}��fiXg�5��ؤ����%��v����=v�����s�M�ő�%�j'B8��K���~^��L�v�u���N��G��vT���q0�|%|�q�\��T�=����X��4Y�U~�
1�9��U��X�7�KBa��:�DM�<�5!AM6|��s�j���b�~aKW�:Sz�5�6�,�G�L/�9�����0�:&��b�9�G�d�4�vm<�h�"S�s�Tf�#�~a�Њm�O����09��BS��H���U��MW�;�_�Vl���Z�c�6W���!�AP���ƭ����=g�#LQa�P,��m�tGa��{��=�	v��r�� I��E�4׽�z.�ʱsyO�GΤ�ĄH�huA��W`���V�;�CꆷD
	?�A�Ka����^Y,]5Z�N	D��e���aZ����e ,Y�u������$c����&����K2���M+��)�]��bh�-�]6�=�WP�L��B0o�}}�}8���*���iz,������c֫�'�)u��v%��
��&j���כ ��r����?G\X�K��@9T��Ix���m5P�y_������T4�;X�
�uZ�,n��_lC�yE*�\�kI7��df��0�����N<�S�ņ�#P�C�qL�k��;\(^R2	�{ݪ��/��Zd	��k��v
�t��:\�x~�H;u<c��c�5Q���]R�n�3��p���ˮ4e�Q�M"W1γ�x��P��c��	ɚ�$wrq�<���h	��7¨[*Ȣ�3�ё��T� �qh�U��03^�:�yV��8����q�BKl&$����No-y8���m�٨��!pD/tD	� nk��?�Jh�����O=/#G�y�c+����Gy��v���Y���~o�R;���5��Ť(t�ڻAw��c~�ؘ]�*L�����^r�0�x�f�q�b�		���X�+z~�w�~;|4V�rEeߞjz��]�Q:��a��,�����\��u�Y��kX�W��O�}CV>l�f"Zee�:���s23������գjE�h��D��l���؍�a�VV���;��yb�A�|�^���	�6o�5��F0��rO�O�xY�w�-�����,
[i�F��EY�Z��G��r�_jb�ԟq��l:&�������t������>s>�'���d,h���`���ğ���fh�\��"���=kP���9ϕA|6�ŀ��W����U��5�%�?��� �2�k%8��[0!��9�o�1�(]�w2�,ݸ����ن�1����g�/��n�mUJ���}�А�
;��>��_.v������BD:�)��l��	+��F�3�]}P�5^�<����U��E��^���[S^��)O��l��!�c"Z@Z&���*���(�����F`_�D���L��i�0Jh������f'C��~�A$��f���>x;-,�c��+�F��&���  5S).Z(%����]�5�nq�VY�A�����V:S��u/'��M?���F������P@'^���If��a��g��Ư�h:N���a%�b:�t{�����˝|� ���t��a�pD��z�ؓ�܏J�F[�oA�QH�B���n�#t0WRw;d�1�b��P�r4�0���U]���+�$��;:�.�ysOJǁ
Zv��r�g�
m��+2?��x�/'�� ��r��A�Ϲ��G�G��+Ȫ~�o���W��$/$'Pi��[w��$�����z��oy�3B�S�I�+
��7�s] ��23e�HE�oC"BtN��lH����'�"<s Y�?�T���_�%k�ʅLQB�R�F8`Ɇ��`������Q����,�g�jNʭ�t�胠T_vo���Y��h��	s|���Ť�$���!��ٻQ2�ɢ�O �jk��'A_����xx���\L�lΛ�
�}���D�|����t��	s��)����a�{�q����IM8�xkk��z[���bH��U����@5'� 7]hK%�m����_���ӷ�눠����q���?tV���.c�[Yp��}�-���AA���L�N��Kb+���!�Π!�}�����Υ.S�l�z��bu�7F{�"*՗KMe�m�~~'�����5;����ZȤx �<��v����M)�ޔQ¥,�M���MY���6�\����ݤ�2�E*�\
�VL��x��t�$�ͬ7R�45aPg1!%�8��0�M _(�"�`,0Nt�p9~D.&�["A�tg3d2�f&^�K+��OJ�;q�l����2\�>�G�0��[Τ!�t�5��6�1��<���]�!p�<��y����#A?3�V������6<I��ǥŒ3�/���@v<��~x�[?����C��Q����]�F��+T7p�|����v:�(~/W�=�Tyd�&����jZ�V)r8\�挙v0	��{����S�����t8t�p���,B��p8S��AFM��b����N�E�����UEi�mt�,?l��O���z#�3�m��	�u��������'(.7�(D�z-Bya�'��d���V��1�~bq���ק������[c)�(�B;�����t�;�ʊV�F$θ;��Y�>ի�MоBl}և��;ߔS�B�d9k���s�� :����1�XC~��Cc��`�bu:�X�_C"�F�D����^/����i��4S� ���s���#DwI���1�����`ʖ3iG~�.��DV��JJ�持j�6�[���OE��i%�:�|�`Ţg���J����!�S�f���O�x1X���OV��ӵε�x]s��!�c�L,hA����F�������2�f���6�8��Y��.##���Qem>3����RU����������LU�P7�kaБƋ(���z�/�o�a~��P�B���0�c�v<7|38P�x�f	�*��	e�;�d=��&o��������t�:��-�-P�0B����N��e��BdPD��p�6�ׂw�/��O�1Ys*]��Q��z\c���&���a�t�b
� �(�)[�����n#x E8�����"��_����M-�"�)�Ψ�)�	D�j'�p\���#u� a�	2������&��O}�Љ0���JLԫg�����}Gg��#íF&�J+A�#���x��0E:~sw��ɧ7ۿ��e�/���uI �c�[Lb92�Q�[2鸌p�Jr�����w��l���o\fh�M�@���w(�����x�Ԕ���=��kL�q춰����;��ؕ���V��i�3Kτ��b0z��XN�hZ,���d�8sfSm����9�,�JԆ�ԍ8������{�t�ؼU��ڔv�v�t~�>�_,m�7w��I�JU�u����э�{TY�X�[_Z�4w���܋8YF��Ym���C�nEjU2���k�6$��B�=]�z�1�8E9�B���c�����In|B��>��g|���s�+g�^�p {�è���E�e��Еe4[z�ĄM�ܐ�,�@��w�Q��E_��e�V]Ĉ��ev틜�*6��t���moLu��։V�!*�=wO�
�����{;+0�woF�Y[|�If�\!ԓ:�判��+K�	@~l��?^�j�D�NM�R����a�Ezw��|:��h�@��X���/^�1��Ozc�����`�oC|���@��v��0B^�4� ��8pR��!4vy��h��j9\�f�^W���\��Y����a�V5���'G�����3��!X���àC�h�s����Wa6a�c��]�6�DB�/��u��Eȿ�!Z��s����(�1�p�� ]����+�,;������m��D�����RM��H�o������Q�B�ו98�?����b��h��!���25s
8�qAJ�O:��*����U��Б�4����
�o�i�Cn�A�
�J��]|��p��6� C�-GL�vs����{s�Q��M�X�tW�i��X_�����)v��d�Xع��w��K=�O�G�6즔�W@��6���z����M�p�xg/�3'n���I�*�'G���K���`|`�&͋)bk'��>c�RD�����h�D�G,7��k�6�����/����Y�'DȤ��.U����ߢ?*�G����n2�o;�!j#��'��H	ۺs����g��f�o$�d;��ͤ�W.����Q�X�1��6d�
�1�8��T^(�*L�?�)	�m��v������S÷�Lo[�_�gN���k��e�y�	�E�̖߅�H�/k���{���_/_�Pa�L�Bo���'�WJ�!{\#i���B�,��fi�N����M��G��0phg�J�Z��&�a�,��gL�T���^�wd�4��fMVb�������sZ:���z��a�*+��(v3,�4�NWuX<&<E�u�?��YݷQ�z͙[�i�d�����W�9g�j�i�N�6��7
M�/��P/,M3!�_��������|�9+�ơ�|�`���(���>Y[�^�z�張A��Mȿ���a���$�n��V�L8�T�yH�QNo��

`(��8�,^O�m�L��������AY���;�a!����Qr�!6|���5as�ԏJ/M��e��UE'1�9X���v�����i��ٛC�g���\3dvj�k�C?:"����A������J8�:{��7��I��8P��sc�Ά#�
�4���� @Ka���F	����~���Ɍڑ2H4M-�g1a�W� x��+�Y��=P��ݴ:F�������^T���~y��P,�;�D�U�*�?no��f�I�Pm�U. tXc���S�>D僰B���� 4q��m���z�v__*��ך�H��ql�7y����X�03�P`2o5��]@�AV�A،$ҡ4X��哟���ze^*����1;���;��a�>F.@�a-�d�������**9�2�,��l�O��U��d�qo&�pQ���̠qG��D�*�O9��'E���)��H��<�۸
�oZ��I�l@��ٚ�JLdd`�kP����æpz&tQJ���W���ˌ�5a���fl�+���T.Q<o�P��p3�w�$v٢h�<`g�,��E���v0T�5��3aw��0�
t�ɰ�C�H������,�@�_��~���d}kѭ#	<�.\q<$~A�A|���gH�:B��aG�;y����[�^��B���1��c� ;`�+ͨ.�$>c2`��O�B0L�.(�kfY#�����x�eH�����U`9�)�G:Xr����F�9g��Kq��MbI�z�X��]�)�@E6���C�8����khQ��nh��BVO>@��+!Z8ɗC-̝���F�_27]Ft
,�r&���׫����R>�=2��*j��Mw�e>�4G=
�s�RE|�G�6���,�(IZ�B\+}�<L���>��f%~>d�sLe{]�R������|p�2�jDl��E�#i�e>��*�B~�Q�&Zک��Z�����j9n����t�;fF��d�y���R���?,���@��(�Xe����~�¥s��(z&�i;�͡/��	����ҧ��glѵ�d��lp�-��z���1Z� ��v���ޟ`,e/3G��X}�G�~�iܟ,����5��2RȬC��M�ᅸ&J�^W%Eu��-Ad�rJҕY,�'��ӫ!����zP(
�_(�	���m(~)��71�ԫ�Н�2�-]s�,uW���+��J����A�Q�/AE�ȁ"i#_o$��S��S[�R�lV�A��j���(��7�ձ��]��L}���BU�����G����l(���4��N����"/���&mm�`�*&�e^p��L�Oi��5r�>��߳m�So�+K�gUHqC�Q�@a�[��K��#oN��#H��Uf��~���Y�T#ѹپI����.����}om:Ў�h^/%n\���e}+�A�*��s���T|A;ƫ����lⱁ�A2��s�v��ͦ�V2�}�l�ֹkg��A�C��0a H��D:_Vԧ b���;�̈PD�7��ئ��Ƈg��j��L����Ut5�-����w��W��u-���MwS�s�����_��U8�*�>3X��l�CP@�j�G/���P��u*���9�p���[�W���L�y�NY�5I,����b/��B�B��T���T`���c�[9{��d�`]t��o�<2=WFt��/U�����b�ƏS��JI(Y��q)au<�t3WEc˭��.*LN���gw����8}�s۪�P�(����]^C��R��Z���׶ �'p:j�TuAL�;��7���13sM�j=P�}A�@$}l��k��玊��O���y{��`�n�6S{^�Ղ�s�b���=؝�����7��_ yݒb��y��Vy��f&���uR��زcz}��LZK�*�����^z�䰖��
̒Sh��y@[��]燢�FT�Vkg�I*
!�C��H�)��|��`S����-A�i�����3�{�xx=��}0�8[p]��"ؑMt��@PUَ:�Q\,�>G����|�Ơ-Gn']F�u_�~��n)qWVaZ��Z�:���Y,m��jܦ4�"��|�Mm�,f'O���߿V���E�*������37��J�<�R��<)��=s���yE�]㸽�r�4��%ؔ����$n��E�${��r��"V&n��kG�t����X��ϙ޴ڛ���j�ф6�O�!�xym(Κ?�]���Xp��DxMs)��(�ڀ���^X�n�q���o++<�w����!���a��iBY�g��V sxڬ���k�(�C�.ˈw�#v$y�ׄr��2
3���ۖ��{��aI��p�+�mr[϶�կ?�����wt��t�#��X�-~���5$3+�@���?^��a�8R]O�3d�����0�aN�B6\�t!'sb
ٳ?F�K�m@����t��&5hي(Hv�8D�_* ���6����;v\�v-L�O$@��k�B����]�Ī\�lG�[U	uK.Xy�.��EI��a�Ҍ��0,~�x��Y�Jk��	LJ�ET�__��aj�XT��Z���2�e>e�He��-����O}$"�@��دM�ʔ�;t��8p���QL�9bݴ�Y���"��D%�����;��Bq�2N!�v�U\��U�ݰ�v�?u����������AM�b�yL�òx�C�X�X� [N)~V� îBĉiN�Z��%�u�hv0w�K��^$qL���hRoA�&6�e��g��6��j�MHv��\��`�K�#�����0�s5N{�U�B�2^"my�;���6��-%���o�fk}	��lMO�_Y�Fޫ�[�!����k38ԩ�H������ �������@x`~,J�o��`�����1��iF8Y�E�";Nǃ�ի֔�>,�Ɍ���J������bVs��lq��PL1||���	��H�kQA�>S��~pt�\�j�x�t1���3κX�Ҟ2,�x�e���ph��zym_��MV��F���F��9-~�#�D����sE*���}݇>�LG�IQ<�k�B�=e�E
�DŢ�����iČ��qc�����"h��1��Ǡ��Nx�=bU��q!̩
 ^?a	��A��R�M/Fl||h|Q�f���g��L;���He*���5�ܲ��L,����T����>o��Ȉ�����UQd
H\�Q�����Ԃ�=�.�L��74H�"�=�ij+����I�!�8W���$8��b.���{	(I��g��}!� CE��̇�ݪ2���Ui�!���Lm0��4ٝ��)�x�Z�=�X+����j������y/򵋍��Y�Y��26�M�Wa���=�� �<=��L����ʂ�g}�br�j��Ɍ*�3�Gs.L2�z8����l@��\���[n�y�Q�7g�*�����3�Os���N�N6�h'}<��,O$���	�d�����.�Lb#�Z&hΑ�ˉoN��L�30����R��ˬQ�BVj6�*z���F��
�"��Q���\��[�d��� .� Aǲ�KJ���g�K�v��1Z��O��h���Z�Lq����H_���o�Я=�N5�6����](�xH@![9#ơ�0��0�i��	�6��Bx-�A�gO�t@� pWZmM�4n��<TW���͵6��#m�䚇�L��)w�'o:�eȈP��wD
��JW PFW��SR^}D[�=�X��۾���K�;.9T�]b#M���̩I��K_�"o"��9%���mf�f�z�M]L��w�XQok���B�!ԢC]��I��*��׹r�0�;�X��k�b�w,��/	��Z6��F�9�#�9.H��2�t�B��1_7U�Zf�5:��a	껤M��G���D	�mp����W����Qm�J�^|��b+X���g��8���h�\���A&?���T��<C�ĭ.�Sa,�p3�9[TcdW�Z���f��m������bqk�����x"�Db��h�Z"f�P��R`�6���q�p�V��� C����ȸ�_�������r9�)cLM��#�N����]BlR���U��(�x�t�n؊��oԅ��q��\ZΚ^D���?"�$ (A�QOz���y���|�3�G<a^X���;�J�\�q.��Vg��)��ѹA{��`�eAYg��Y��#��w�lPi*�m[����h�Ħv4����P����s�a=�ݵ����h�5��Ԩ0���m�h�y��6���(v����
)�G�`4�|vx�S�R��.�����`��,�#J�E5O���b��!��f��G��u����H˽
ƨgzԪ�ؙ;��R(R����E����v�9&��Zi�;[����!2�xǛ-����;͔/8-�����4��c��"�k�S@�Y֏��7l��<Z��M��;�/�G��~f��{��&�C�n�!�OF!|�+�˅���sk3R��çm ����֍�RY��D>���l��3=@~�3'�(�,h�7C£���?_��Gt/�ϰ�la���J�7�J"(R�x���PwP$F�Ͱ��+!�;���֑����.�l=5̽|�wd�%���:��c�C�6�=��7]��M�ppt�_��k}�:��̯�u�a=c�.�~b���B���2/��:�6�<pp-"�y����D;�5��+���L��V��؅2 ��"/����S��{2���b�U�3�S��L����g��8Z(���-(�E�ٌ����8�v�'��R�7�wߊH��l�m`��f�s?^1J/�GS���CAtVy��t^K)F��eW~3����7��>���f�B�딓��ÿ�9o�����6�Z�z�Q��X.Z�[�xaUW��ǫ��1���u�s�d~��^}�3��sN�0*9��2����,'Kd,�MYyBY{���=�zDn�|I��򢔯3c��ja���gť���V�Yu.�m��F�;�qq<u+@@���KW	��M������a�q���I�m��)�q'4���=�Үǅ ]4���#��&OG1Ix�(����i�]=��'��2���8���,���GÆ���Q�+|�-�9f�ɩ����GGB4��?�E���k�5ɭ�X#��۵?��n�����jT��j�w����"��|�*5�uK���d�}���x���d�r�oB|��/��ha,���}9�����s����F#����
���Tb�mTV���B`mX.��Y�ϐC[.�b�.K�-}�no�B?�9���W�J9hj�&|�����m̺�m⌑���y�fS�1�{ͤ�<v�\.t���O3����u(�%/T!)D��!��e�Zz����
�n?'�r�(X^Q�[��ʡ�O��42x�#��=o�z��Ն>#E��[���W���JY�%��]oy�"��(Dvqopa�p��׹w�?7������P
˙%"�D��s��}���"���:v5���`��tAU����ɖG~t�/�w)HSY%�Bb7K��y�'Ch"s��il�� �nˋ�2�Z�e�W�"�����>s�|�v��ӄ����61J~{���0���4B���"�M�J���:ut"k9\SPnH[&0v�9�!����s��OpN� ��bN��B^X}��٠d��z�xYs����Q|�N��
p���s٪w�EV��r+�)��>�]O�����L�v�� ���(�c]� ���@�������ὀD�ձ���˸�������
�{s5=ܺH��q*�t#x�M�*8�[�v}�$���H�j�~�˶v�� ��Z�'�B�oJ0��\g���;X�����:��mjz	4�o!T�xe�Cr���ps�_s�#�]$�>�J��*�a[���}���z��Rt��P:e�:��J;���z���lmH =�`Oܮ�c���X�^\����sX�V���X��q������B`��5P��p�C�Bۧr�׈����٪Y��7Z�制�y0��+z� Y�[f�~+�Ӎ"��I����w58��*��+��8�@��3In��U����d��X@o�ᇤ����C��X����Ę3rIi+��|�??�����b<�m�!����Z���d~�U������F5�)Fڽ�Gp�/J��[u�	ve;k��6�~��P�
��C"��If��\�A?�ө��u���s\ۅ�zy]+��XH��9��3K?>�]�&M1a�6Q`������f��F�\��H�N��z�[�2ԝp�8�/C~V���9ԩ��yOZT�@�=���@�óf)�cL��&��# C*9Wó�y�А�L�O�u���j��4V�n�'��z*;<��/,�6ὔ����f�Qܖ��b�h߸pry�e�Tz*Z��i������ւ����AǙ�X�����h?�i<!i�p��j�	�C����3�5x���zq����=���è?)D�r҆M��-�kO����^�B�F�5�|�e
6!3�ץ�g�|ݏI�޹��#ZW�?��Ċ�������^��r�����Q�Ґ8��ML��p�G�nC8 �4�gg�N�����M�c��G�\i1P�s�pS�g�WJ'"l44�m^�rzT/����|"�3}(���*�@��skFE�A�`�0��$�F�U��m�*EZ	�n���{n9 6��A<~\���:$>�3��29����[�aH�_�u9�Ё}���?���[�	���aS�k�qˣ�ZK+Dړ,H�{����Q�tS�IQ?�=�Yn���*��Ԁ�^z*~��c�Y,M���ZD���.�7V)����0�SCi�S�&�Y�i��t p�ÞD�yz�|l���x������S@�.��\2�m7jA�~8S3�#R��Lݒ����y�f���e�Z���UU�j�+�VС�X��Ǣ��J/����x��{�A�
�&]�ZPc�#`N�6���f��0�����8P`%O�n���*�����9l�bR�q�y&uǅwyɼ���ź�AӘg"�5Z�'��ƿK�N�mY#��%yQ�R	+�ng��v�l�����)����Tws?x�f��ǉjrI=m$ؾ�]tX;���^��A������E9&�|v��z �}��'u>pn!�B���$7sL�����ے/J��)��"�k�R�
��� �����E>�r�g�dp��DqdY3����<�%ȓo	U�!$'�"��9�`.FXl'S��(N��d�"MyJ:ܐ]D=�_��G�q\�ߐ�:�t ���m�̀�4�7��9�G��l@�������.�n˖�Ǥ?�U�E*3��2+E���x��-�JS��`��051q~ɍ�'�3`m�F�Ó�2
E��|$w�T�'��D�j��\{�(��a�5<]�/b.(��`*v�|Fw�vo��=��9'w�R|��S�{�y��ұCJ�N�d�x�Xo��1"�ʠ��e`�n��`��ӡ��'���3�\�i��c���ƪ��X��햠�C�W���K-��n���,z�ƌl%��߫ ��Z-�@�̖qh��1�6��#ݧnKQ���HX�R�h�a�R�w8���I�j����C�)o4\�I�{-�MZQߐ0A5���YO�������x͍ ���.*��ί%��OSA Jcj����`N�\��oS$����&'� b���l��?�;c����^~1x��D�28d���}�[4C��tޞ{������zJ���8�TX'�����!�ËwR:C���5�'wf5�b���Ո"���z��.բl7��x����j�
� �T{�n f40���	�h�㛓��~gy&��xA�F�PwH���>eO��eV�mM��^�b%����/C,#=2�CQ#����iŐD��X��v��o�g|E�ɷ|��W��R���͕}�k��ԝL���3�34�y�'o�8�S�)z��&���U���r�D"��v*>�D�DP�Î����,	D;-���L��0�oG�郒
5 '`��`�A�v%Fi�6�n��5�`�s�0C7����VƯ�Jm'~��vw�])p�Z��S�hn�D']�ЫDX�)�I�$|Vu��g8
T�xˮ�J8�C�O��b���Y����% 1b%�`*il�\U��u1�2[;���H�oN�e��ɯ���z��ۡ�ɿ퓽,�~����m�O�$�qͫ�J8�<b����G|vܨz�HQՒH���Ir�j0��W�<{ZwWkN�R�qa���]]!sӧmv0 �t�B�҄�S��*�]Ϥ��I����{kY�ص�v
���5�KD��R:u����*gȾ�gG�ӗ�����鵻�Ə}2�ȇl`������](�z�[�}K��Fq][���),���̋�E�\Vp7�8~�ꑐ;:`���T$Op�od:���jF�T�������+?�Q{�!�"���dAcTw73<,$ S�i�����v	v��-����r�dm����k�#�ylfV*��3�$D��Q�|��+�Y��|���r�}���\_��xhk�h�[� 7b
�Xk����@l,��~9f�̟�Jgb�ФF�R��Iŏ2$$�ѧ��p��OOJq�����$��ꦷ��@�x�.~����)���yݺ.��x y�H<j�g�&ΖK.�g�_�Hd���s�=��Vq�.�N����D�h���?���T�~�oDa�S�yt�r�r��8$�;p�#��?	���b
�#��Q҃���Z��\uh��p�2��F����!Y�-�R�v���ڡ�"1	b�@�����D��,���z���Q��/U��'�Du�\��P�0���X�����2=���y����X
��ߵIoO�2|�K��"�V�m����튺�BU�qNEg��}/]�7����L�?��Gh�!\Ǟ�~�ėC��A���o#�t@H��D��7���aʆ��;�UR���� k���[������mq��<�w~G�����^5�����~!��9m)hɭ�����1q��s���K]�v>N�������-�I[��p��UrBI��$0�էy�L�2��:e�G�T�(*>�{��p��֎�3Ո�F(y�͙΍7�5_�e�0�Grlh��N�4���y}sx� KJd�@b	��:�~���U��w��OgQ`�(�����3ǀ" -�xģ�A��9ŴƔ?�%���� {ѵgD>������ �,�A6y{Yy�ݭ��'ND�	�x����H햧v���MP��ݤ8�-���~ k�a�_�
�")���K�"��g^ya�`�3tb�f���"��B"�H3�> s�_��-����s�빂�=����]k�E�����O�א�͌,Yn�R'ͥ�Sx��Ί��F��-��d�L� N�q	&�>�%x�V���2�2��>�b�ۘ/��