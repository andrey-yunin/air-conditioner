-- embedded_computer_system.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity embedded_computer_system is
	port (
		clk_clk                        : in    std_logic                     := '0';             --                    clk.clk
		pio_0_export                   : out   std_logic_vector(7 downto 0);                     --                  pio_0.export
		pll_c1_clk                     : out   std_logic;                                        --                 pll_c1.clk
		reset_reset_n                  : in    std_logic                     := '0';             --                  reset.reset_n
		sdram_controller_addr          : out   std_logic_vector(12 downto 0);                    --       sdram_controller.addr
		sdram_controller_ba            : out   std_logic_vector(1 downto 0);                     --                       .ba
		sdram_controller_cas_n         : out   std_logic;                                        --                       .cas_n
		sdram_controller_cke           : out   std_logic;                                        --                       .cke
		sdram_controller_cs_n          : out   std_logic;                                        --                       .cs_n
		sdram_controller_dq            : inout std_logic_vector(15 downto 0) := (others => '0'); --                       .dq
		sdram_controller_dqm           : out   std_logic_vector(1 downto 0);                     --                       .dqm
		sdram_controller_ras_n         : out   std_logic;                                        --                       .ras_n
		sdram_controller_we_n          : out   std_logic;                                        --                       .we_n
		sierra_0_conduit_end_export    : out   std_logic_vector(2 downto 0);                     --   sierra_0_conduit_end.export
		sierra_0_conduit_end_1_export  : in    std_logic_vector(1 downto 0)  := (others => '0'); -- sierra_0_conduit_end_1.export
		temperature_set_ip_0_writedata : in    std_logic_vector(1 downto 0)  := (others => '0'); --   temperature_set_ip_0.writedata
		vga_ip_0_conduit_end_vga_b     : out   std_logic_vector(3 downto 0);                     --   vga_ip_0_conduit_end.vga_b
		vga_ip_0_conduit_end_vga_g     : out   std_logic_vector(3 downto 0);                     --                       .vga_g
		vga_ip_0_conduit_end_vga_r     : out   std_logic_vector(3 downto 0);                     --                       .vga_r
		vga_ip_0_conduit_end_vga_vs    : out   std_logic;                                        --                       .vga_vs
		vga_ip_0_conduit_end_vga_hs    : out   std_logic                                         --                       .vga_hs
	);
end entity embedded_computer_system;

architecture rtl of embedded_computer_system is
	component VGA_IP is
		port (
			data_controller_in    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			wren_controller       : in  std_logic                     := 'X';             -- write
			cs_n                  : in  std_logic                     := 'X';             -- chipselect_n
			address_controller_in : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			reset_controller      : in  std_logic                     := 'X';             -- reset_n
			CLOCK_controller_50   : in  std_logic                     := 'X';             -- clk
			VGA_controller_B      : out std_logic_vector(3 downto 0);                     -- vga_b
			VGA_controller_G      : out std_logic_vector(3 downto 0);                     -- vga_g
			VGA_controller_R      : out std_logic_vector(3 downto 0);                     -- vga_r
			VGA_controller_VS     : out std_logic;                                        -- vga_vs
			VGA_controller_HS     : out std_logic                                         -- vga_hs
		);
	end component VGA_IP;

	component embedded_computer_system_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component embedded_computer_system_cpu;

	component embedded_computer_system_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component embedded_computer_system_jtag_uart;

	component embedded_computer_system_modular_adc_0 is
		generic (
			is_this_first_or_second_adc : integer := 1
		);
		port (
			clock_clk                  : in  std_logic                     := 'X';             -- clk
			reset_sink_reset_n         : in  std_logic                     := 'X';             -- reset_n
			adc_pll_clock_clk          : in  std_logic                     := 'X';             -- clk
			adc_pll_locked_export      : in  std_logic                     := 'X';             -- export
			sequencer_csr_address      : in  std_logic                     := 'X';             -- address
			sequencer_csr_read         : in  std_logic                     := 'X';             -- read
			sequencer_csr_write        : in  std_logic                     := 'X';             -- write
			sequencer_csr_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sequencer_csr_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			sample_store_csr_address   : in  std_logic_vector(6 downto 0)  := (others => 'X'); -- address
			sample_store_csr_read      : in  std_logic                     := 'X';             -- read
			sample_store_csr_write     : in  std_logic                     := 'X';             -- write
			sample_store_csr_writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			sample_store_csr_readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			sample_store_irq_irq       : out std_logic                                         -- irq
		);
	end component embedded_computer_system_modular_adc_0;

	component embedded_computer_system_pio_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component embedded_computer_system_pio_0;

	component embedded_computer_system_pll is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			c2                 : out std_logic;                                        -- clk
			locked             : out std_logic;                                        -- export
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component embedded_computer_system_pll;

	component embedded_computer_system_sdram_controller is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component embedded_computer_system_sdram_controller;

	component sierra is
		port (
			address                     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			chipselect_n                : in  std_logic                     := 'X';             -- chipselect_n
			read_n                      : in  std_logic                     := 'X';             -- read_n
			writedata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			write_n                     : in  std_logic                     := 'X';             -- write_n
			readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			clk                         : in  std_logic                     := 'X';             -- clk
			reset_n                     : in  std_logic                     := 'X';             -- reset_n
			external_runing_taskid_info : out std_logic_vector(2 downto 0);                     -- export
			irq                         : out std_logic;                                        -- irq
			extirq_n                    : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component sierra;

	component embedded_computer_system_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component embedded_computer_system_sysid_qsys_0;

	component temperature_set_IP is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			cs_n     : in  std_logic                     := 'X';             -- chipselect_n
			read_n   : in  std_logic                     := 'X';             -- read_n
			data_out : out std_logic_vector(31 downto 0);                    -- readdata
			data_in  : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- writedata
		);
	end component temperature_set_IP;

	component embedded_computer_system_value_0 is
		port (
			avs_a_read         : in  std_logic                     := 'X';             -- read
			avs_a_write        : in  std_logic                     := 'X';             -- write
			avs_a_address      : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			avs_a_writedata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avs_a_byteenable   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avs_a_readdata     : out std_logic_vector(31 downto 0);                    -- readdata
			avs_cra_read       : in  std_logic                     := 'X';             -- read
			avs_cra_write      : in  std_logic                     := 'X';             -- write
			avs_cra_address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			avs_cra_writedata  : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			avs_cra_byteenable : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			avs_cra_readdata   : out std_logic_vector(63 downto 0);                    -- readdata
			clock              : in  std_logic                     := 'X';             -- clk
			done_irq           : out std_logic;                                        -- irq
			resetn             : in  std_logic                     := 'X'              -- reset_n
		);
	end component embedded_computer_system_value_0;

	component embedded_computer_system_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                         : in  std_logic                     := 'X';             -- clk
			pll_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset                 : in  std_logic                     := 'X';             -- reset
			jtag_uart_reset_reset_bridge_in_reset_reset           : in  std_logic                     := 'X';             -- reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                               : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                           : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                  : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                              : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                                 : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                           : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                        : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                    : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                           : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_debug_mem_slave_address                           : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                             : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                              : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess                       : out std_logic;                                        -- debugaccess
			jtag_uart_avalon_jtag_slave_address                   : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                     : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                      : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                : out std_logic;                                        -- chipselect
			modular_adc_0_sample_store_csr_address                : out std_logic_vector(6 downto 0);                     -- address
			modular_adc_0_sample_store_csr_write                  : out std_logic;                                        -- write
			modular_adc_0_sample_store_csr_read                   : out std_logic;                                        -- read
			modular_adc_0_sample_store_csr_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			modular_adc_0_sample_store_csr_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			modular_adc_0_sequencer_csr_address                   : out std_logic_vector(0 downto 0);                     -- address
			modular_adc_0_sequencer_csr_write                     : out std_logic;                                        -- write
			modular_adc_0_sequencer_csr_read                      : out std_logic;                                        -- read
			modular_adc_0_sequencer_csr_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			modular_adc_0_sequencer_csr_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			pio_0_s1_address                                      : out std_logic_vector(1 downto 0);                     -- address
			pio_0_s1_write                                        : out std_logic;                                        -- write
			pio_0_s1_readdata                                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_0_s1_writedata                                    : out std_logic_vector(31 downto 0);                    -- writedata
			pio_0_s1_chipselect                                   : out std_logic;                                        -- chipselect
			pll_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pll_pll_slave_write                                   : out std_logic;                                        -- write
			pll_pll_slave_read                                    : out std_logic;                                        -- read
			pll_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			sdram_controller_s1_address                           : out std_logic_vector(24 downto 0);                    -- address
			sdram_controller_s1_write                             : out std_logic;                                        -- write
			sdram_controller_s1_read                              : out std_logic;                                        -- read
			sdram_controller_s1_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_controller_s1_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_controller_s1_byteenable                        : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_controller_s1_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			sdram_controller_s1_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			sdram_controller_s1_chipselect                        : out std_logic;                                        -- chipselect
			sierra_0_avalon_slave_0_address                       : out std_logic_vector(7 downto 0);                     -- address
			sierra_0_avalon_slave_0_write                         : out std_logic;                                        -- write
			sierra_0_avalon_slave_0_read                          : out std_logic;                                        -- read
			sierra_0_avalon_slave_0_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sierra_0_avalon_slave_0_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			sierra_0_avalon_slave_0_chipselect                    : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address                    : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			temperature_set_IP_0_avalon_slave_0_read              : out std_logic;                                        -- read
			temperature_set_IP_0_avalon_slave_0_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			temperature_set_IP_0_avalon_slave_0_chipselect        : out std_logic;                                        -- chipselect
			value_0_avs_a_address                                 : out std_logic_vector(5 downto 0);                     -- address
			value_0_avs_a_write                                   : out std_logic;                                        -- write
			value_0_avs_a_read                                    : out std_logic;                                        -- read
			value_0_avs_a_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			value_0_avs_a_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			value_0_avs_a_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			value_0_avs_cra_address                               : out std_logic_vector(2 downto 0);                     -- address
			value_0_avs_cra_write                                 : out std_logic;                                        -- write
			value_0_avs_cra_read                                  : out std_logic;                                        -- read
			value_0_avs_cra_readdata                              : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			value_0_avs_cra_writedata                             : out std_logic_vector(63 downto 0);                    -- writedata
			value_0_avs_cra_byteenable                            : out std_logic_vector(7 downto 0);                     -- byteenable
			VGA_IP_0_avalon_slave_0_address                       : out std_logic_vector(16 downto 0);                    -- address
			VGA_IP_0_avalon_slave_0_write                         : out std_logic;                                        -- write
			VGA_IP_0_avalon_slave_0_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			VGA_IP_0_avalon_slave_0_chipselect                    : out std_logic                                         -- chipselect
		);
	end component embedded_computer_system_mm_interconnect_0;

	component embedded_computer_system_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component embedded_computer_system_irq_mapper;

	component embedded_computer_system_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component embedded_computer_system_rst_controller;

	component embedded_computer_system_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component embedded_computer_system_rst_controller_001;

	signal pll_c0_clk                                                                 : std_logic;                     -- pll:c0 -> [VGA_IP_0:CLOCK_controller_50, cpu:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:pll_c0_clk, modular_adc_0:clock_clk, pio_0:clk, rst_controller:clk, rst_controller_001:clk, sdram_controller:clk, sierra_0:clk, sysid_qsys_0:clock, temperature_set_IP_0:clk, value_0:clock]
	signal pll_c2_clk                                                                 : std_logic;                     -- pll:c2 -> modular_adc_0:adc_pll_clock_clk
	signal pll_locked_conduit_export                                                  : std_logic;                     -- pll:locked -> modular_adc_0:adc_pll_locked_export
	signal cpu_data_master_readdata                                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                                : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                                : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                                    : std_logic_vector(27 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                                 : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                                       : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                                      : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                                  : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                         : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                             : std_logic_vector(27 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                                : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect                   : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata                     : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest                  : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address                      : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                         : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                        : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect                       : std_logic;                     -- mm_interconnect_0:VGA_IP_0_avalon_slave_0_chipselect -> mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect:in
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_address                          : std_logic_vector(16 downto 0); -- mm_interconnect_0:VGA_IP_0_avalon_slave_0_address -> VGA_IP_0:address_controller_in
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_write                            : std_logic;                     -- mm_interconnect_0:VGA_IP_0_avalon_slave_0_write -> VGA_IP_0:wren_controller
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:VGA_IP_0_avalon_slave_0_writedata -> VGA_IP_0:data_controller_in
	signal mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_chipselect           : std_logic;                     -- mm_interconnect_0:temperature_set_IP_0_avalon_slave_0_chipselect -> mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_chipselect:in
	signal mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_readdata             : std_logic_vector(31 downto 0); -- temperature_set_IP_0:data_out -> mm_interconnect_0:temperature_set_IP_0_avalon_slave_0_readdata
	signal mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_read                 : std_logic;                     -- mm_interconnect_0:temperature_set_IP_0_avalon_slave_0_read -> mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_read:in
	signal mm_interconnect_0_sierra_0_avalon_slave_0_chipselect                       : std_logic;                     -- mm_interconnect_0:sierra_0_avalon_slave_0_chipselect -> mm_interconnect_0_sierra_0_avalon_slave_0_chipselect:in
	signal mm_interconnect_0_sierra_0_avalon_slave_0_readdata                         : std_logic_vector(31 downto 0); -- sierra_0:readdata -> mm_interconnect_0:sierra_0_avalon_slave_0_readdata
	signal mm_interconnect_0_sierra_0_avalon_slave_0_address                          : std_logic_vector(7 downto 0);  -- mm_interconnect_0:sierra_0_avalon_slave_0_address -> sierra_0:address
	signal mm_interconnect_0_sierra_0_avalon_slave_0_read                             : std_logic;                     -- mm_interconnect_0:sierra_0_avalon_slave_0_read -> mm_interconnect_0_sierra_0_avalon_slave_0_read:in
	signal mm_interconnect_0_sierra_0_avalon_slave_0_write                            : std_logic;                     -- mm_interconnect_0:sierra_0_avalon_slave_0_write -> mm_interconnect_0_sierra_0_avalon_slave_0_write:in
	signal mm_interconnect_0_sierra_0_avalon_slave_0_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:sierra_0_avalon_slave_0_writedata -> sierra_0:writedata
	signal mm_interconnect_0_value_0_avs_a_readdata                                   : std_logic_vector(31 downto 0); -- value_0:avs_a_readdata -> mm_interconnect_0:value_0_avs_a_readdata
	signal mm_interconnect_0_value_0_avs_a_address                                    : std_logic_vector(5 downto 0);  -- mm_interconnect_0:value_0_avs_a_address -> value_0:avs_a_address
	signal mm_interconnect_0_value_0_avs_a_read                                       : std_logic;                     -- mm_interconnect_0:value_0_avs_a_read -> value_0:avs_a_read
	signal mm_interconnect_0_value_0_avs_a_byteenable                                 : std_logic_vector(3 downto 0);  -- mm_interconnect_0:value_0_avs_a_byteenable -> value_0:avs_a_byteenable
	signal mm_interconnect_0_value_0_avs_a_write                                      : std_logic;                     -- mm_interconnect_0:value_0_avs_a_write -> value_0:avs_a_write
	signal mm_interconnect_0_value_0_avs_a_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:value_0_avs_a_writedata -> value_0:avs_a_writedata
	signal mm_interconnect_0_value_0_avs_cra_readdata                                 : std_logic_vector(63 downto 0); -- value_0:avs_cra_readdata -> mm_interconnect_0:value_0_avs_cra_readdata
	signal mm_interconnect_0_value_0_avs_cra_address                                  : std_logic_vector(2 downto 0);  -- mm_interconnect_0:value_0_avs_cra_address -> value_0:avs_cra_address
	signal mm_interconnect_0_value_0_avs_cra_read                                     : std_logic;                     -- mm_interconnect_0:value_0_avs_cra_read -> value_0:avs_cra_read
	signal mm_interconnect_0_value_0_avs_cra_byteenable                               : std_logic_vector(7 downto 0);  -- mm_interconnect_0:value_0_avs_cra_byteenable -> value_0:avs_cra_byteenable
	signal mm_interconnect_0_value_0_avs_cra_write                                    : std_logic;                     -- mm_interconnect_0:value_0_avs_cra_write -> value_0:avs_cra_write
	signal mm_interconnect_0_value_0_avs_cra_writedata                                : std_logic_vector(63 downto 0); -- mm_interconnect_0:value_0_avs_cra_writedata -> value_0:avs_cra_writedata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata                      : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address                       : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                             : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                          : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                          : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                              : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                                 : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                                : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_pll_pll_slave_readdata                                   : std_logic_vector(31 downto 0); -- pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	signal mm_interconnect_0_pll_pll_slave_address                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pll_pll_slave_address -> pll:address
	signal mm_interconnect_0_pll_pll_slave_read                                       : std_logic;                     -- mm_interconnect_0:pll_pll_slave_read -> pll:read
	signal mm_interconnect_0_pll_pll_slave_write                                      : std_logic;                     -- mm_interconnect_0:pll_pll_slave_write -> pll:write
	signal mm_interconnect_0_pll_pll_slave_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	signal mm_interconnect_0_sdram_controller_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	signal mm_interconnect_0_sdram_controller_s1_readdata                             : std_logic_vector(15 downto 0); -- sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	signal mm_interconnect_0_sdram_controller_s1_waitrequest                          : std_logic;                     -- sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	signal mm_interconnect_0_sdram_controller_s1_address                              : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	signal mm_interconnect_0_sdram_controller_s1_read                                 : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_read -> mm_interconnect_0_sdram_controller_s1_read:in
	signal mm_interconnect_0_sdram_controller_s1_byteenable                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_controller_s1_byteenable -> mm_interconnect_0_sdram_controller_s1_byteenable:in
	signal mm_interconnect_0_sdram_controller_s1_readdatavalid                        : std_logic;                     -- sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	signal mm_interconnect_0_sdram_controller_s1_write                                : std_logic;                     -- mm_interconnect_0:sdram_controller_s1_write -> mm_interconnect_0_sdram_controller_s1_write:in
	signal mm_interconnect_0_sdram_controller_s1_writedata                            : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	signal mm_interconnect_0_pio_0_s1_chipselect                                      : std_logic;                     -- mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	signal mm_interconnect_0_pio_0_s1_readdata                                        : std_logic_vector(31 downto 0); -- pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	signal mm_interconnect_0_pio_0_s1_address                                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_0_s1_address -> pio_0:address
	signal mm_interconnect_0_pio_0_s1_write                                           : std_logic;                     -- mm_interconnect_0:pio_0_s1_write -> mm_interconnect_0_pio_0_s1_write:in
	signal mm_interconnect_0_pio_0_s1_writedata                                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	signal mm_interconnect_0_modular_adc_0_sample_store_csr_readdata                  : std_logic_vector(31 downto 0); -- modular_adc_0:sample_store_csr_readdata -> mm_interconnect_0:modular_adc_0_sample_store_csr_readdata
	signal mm_interconnect_0_modular_adc_0_sample_store_csr_address                   : std_logic_vector(6 downto 0);  -- mm_interconnect_0:modular_adc_0_sample_store_csr_address -> modular_adc_0:sample_store_csr_address
	signal mm_interconnect_0_modular_adc_0_sample_store_csr_read                      : std_logic;                     -- mm_interconnect_0:modular_adc_0_sample_store_csr_read -> modular_adc_0:sample_store_csr_read
	signal mm_interconnect_0_modular_adc_0_sample_store_csr_write                     : std_logic;                     -- mm_interconnect_0:modular_adc_0_sample_store_csr_write -> modular_adc_0:sample_store_csr_write
	signal mm_interconnect_0_modular_adc_0_sample_store_csr_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:modular_adc_0_sample_store_csr_writedata -> modular_adc_0:sample_store_csr_writedata
	signal mm_interconnect_0_modular_adc_0_sequencer_csr_readdata                     : std_logic_vector(31 downto 0); -- modular_adc_0:sequencer_csr_readdata -> mm_interconnect_0:modular_adc_0_sequencer_csr_readdata
	signal mm_interconnect_0_modular_adc_0_sequencer_csr_address                      : std_logic_vector(0 downto 0);  -- mm_interconnect_0:modular_adc_0_sequencer_csr_address -> modular_adc_0:sequencer_csr_address
	signal mm_interconnect_0_modular_adc_0_sequencer_csr_read                         : std_logic;                     -- mm_interconnect_0:modular_adc_0_sequencer_csr_read -> modular_adc_0:sequencer_csr_read
	signal mm_interconnect_0_modular_adc_0_sequencer_csr_write                        : std_logic;                     -- mm_interconnect_0:modular_adc_0_sequencer_csr_write -> modular_adc_0:sequencer_csr_write
	signal mm_interconnect_0_modular_adc_0_sequencer_csr_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:modular_adc_0_sequencer_csr_writedata -> modular_adc_0:sequencer_csr_writedata
	signal irq_mapper_receiver0_irq                                                   : std_logic;                     -- sierra_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                   : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                   : std_logic;                     -- value_0:done_irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                   : std_logic;                     -- modular_adc_0:sample_store_irq_irq -> irq_mapper:receiver3_irq
	signal cpu_irq_irq                                                                : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                             : std_logic;                     -- rst_controller:reset_out -> [mm_interconnect_0:jtag_uart_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in]
	signal cpu_debug_reset_request_reset                                              : std_logic;                     -- cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_002:reset_in1]
	signal rst_controller_001_reset_out_reset                                         : std_logic;                     -- rst_controller_001:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                                     : std_logic;                     -- rst_controller_001:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	signal rst_controller_002_reset_out_reset                                         : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]
	signal reset_reset_n_ports_inv                                                    : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv               : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv              : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect_ports_inv             : std_logic;                     -- mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect:inv -> VGA_IP_0:cs_n
	signal mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_chipselect_ports_inv : std_logic;                     -- mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_chipselect:inv -> temperature_set_IP_0:cs_n
	signal mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_read_ports_inv       : std_logic;                     -- mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_read:inv -> temperature_set_IP_0:read_n
	signal mm_interconnect_0_sierra_0_avalon_slave_0_chipselect_ports_inv             : std_logic;                     -- mm_interconnect_0_sierra_0_avalon_slave_0_chipselect:inv -> sierra_0:chipselect_n
	signal mm_interconnect_0_sierra_0_avalon_slave_0_read_ports_inv                   : std_logic;                     -- mm_interconnect_0_sierra_0_avalon_slave_0_read:inv -> sierra_0:read_n
	signal mm_interconnect_0_sierra_0_avalon_slave_0_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_sierra_0_avalon_slave_0_write:inv -> sierra_0:write_n
	signal mm_interconnect_0_sdram_controller_s1_read_ports_inv                       : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_read:inv -> sdram_controller:az_rd_n
	signal mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_controller_s1_byteenable:inv -> sdram_controller:az_be_n
	signal mm_interconnect_0_sdram_controller_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_sdram_controller_s1_write:inv -> sdram_controller:az_wr_n
	signal mm_interconnect_0_pio_0_s1_write_ports_inv                                 : std_logic;                     -- mm_interconnect_0_pio_0_s1_write:inv -> pio_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                                   : std_logic;                     -- rst_controller_reset_out_reset:inv -> [VGA_IP_0:reset_controller, jtag_uart:rst_n, modular_adc_0:reset_sink_reset_n, pio_0:reset_n, sdram_controller:reset_n, sysid_qsys_0:reset_n, temperature_set_IP_0:reset_n, value_0:resetn]
	signal rst_controller_001_reset_out_reset_ports_inv                               : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [cpu:reset_n, sierra_0:reset_n]

begin

	vga_ip_0 : component VGA_IP
		port map (
			data_controller_in    => mm_interconnect_0_vga_ip_0_avalon_slave_0_writedata,            -- avalon_slave_0.writedata
			wren_controller       => mm_interconnect_0_vga_ip_0_avalon_slave_0_write,                --               .write
			cs_n                  => mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect_ports_inv, --               .chipselect_n
			address_controller_in => mm_interconnect_0_vga_ip_0_avalon_slave_0_address,              --               .address
			reset_controller      => rst_controller_reset_out_reset_ports_inv,                       --          reset.reset_n
			CLOCK_controller_50   => pll_c0_clk,                                                     --          clock.clk
			VGA_controller_B      => vga_ip_0_conduit_end_vga_b,                                     --    conduit_end.vga_b
			VGA_controller_G      => vga_ip_0_conduit_end_vga_g,                                     --               .vga_g
			VGA_controller_R      => vga_ip_0_conduit_end_vga_r,                                     --               .vga_r
			VGA_controller_VS     => vga_ip_0_conduit_end_vga_vs,                                    --               .vga_vs
			VGA_controller_HS     => vga_ip_0_conduit_end_vga_hs                                     --               .vga_hs
		);

	cpu : component embedded_computer_system_cpu
		port map (
			clk                                 => pll_c0_clk,                                        --                       clk.clk
			reset_n                             => rst_controller_001_reset_out_reset_ports_inv,      --                     reset.reset_n
			reset_req                           => rst_controller_001_reset_out_reset_req,            --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	jtag_uart : component embedded_computer_system_jtag_uart
		port map (
			clk            => pll_c0_clk,                                                    --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	modular_adc_0 : component embedded_computer_system_modular_adc_0
		generic map (
			is_this_first_or_second_adc => 1
		)
		port map (
			clock_clk                  => pll_c0_clk,                                                 --            clock.clk
			reset_sink_reset_n         => rst_controller_reset_out_reset_ports_inv,                   --       reset_sink.reset_n
			adc_pll_clock_clk          => pll_c2_clk,                                                 --    adc_pll_clock.clk
			adc_pll_locked_export      => pll_locked_conduit_export,                                  --   adc_pll_locked.export
			sequencer_csr_address      => mm_interconnect_0_modular_adc_0_sequencer_csr_address(0),   --    sequencer_csr.address
			sequencer_csr_read         => mm_interconnect_0_modular_adc_0_sequencer_csr_read,         --                 .read
			sequencer_csr_write        => mm_interconnect_0_modular_adc_0_sequencer_csr_write,        --                 .write
			sequencer_csr_writedata    => mm_interconnect_0_modular_adc_0_sequencer_csr_writedata,    --                 .writedata
			sequencer_csr_readdata     => mm_interconnect_0_modular_adc_0_sequencer_csr_readdata,     --                 .readdata
			sample_store_csr_address   => mm_interconnect_0_modular_adc_0_sample_store_csr_address,   -- sample_store_csr.address
			sample_store_csr_read      => mm_interconnect_0_modular_adc_0_sample_store_csr_read,      --                 .read
			sample_store_csr_write     => mm_interconnect_0_modular_adc_0_sample_store_csr_write,     --                 .write
			sample_store_csr_writedata => mm_interconnect_0_modular_adc_0_sample_store_csr_writedata, --                 .writedata
			sample_store_csr_readdata  => mm_interconnect_0_modular_adc_0_sample_store_csr_readdata,  --                 .readdata
			sample_store_irq_irq       => irq_mapper_receiver3_irq                                    -- sample_store_irq.irq
		);

	pio_0 : component embedded_computer_system_pio_0
		port map (
			clk        => pll_c0_clk,                                 --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address    => mm_interconnect_0_pio_0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_0_s1_readdata,        --                    .readdata
			out_port   => pio_0_export                                -- external_connection.export
		);

	pll : component embedded_computer_system_pll
		port map (
			clk                => clk_clk,                                   --       inclk_interface.clk
			reset              => rst_controller_002_reset_out_reset,        -- inclk_interface_reset.reset
			read               => mm_interconnect_0_pll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_pll_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_pll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_pll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_pll_pll_slave_writedata, --                      .writedata
			c0                 => pll_c0_clk,                                --                    c0.clk
			c1                 => pll_c1_clk,                                --                    c1.clk
			c2                 => pll_c2_clk,                                --                    c2.clk
			locked             => pll_locked_conduit_export,                 --        locked_conduit.export
			scandone           => open,                                      --           (terminated)
			scandataout        => open,                                      --           (terminated)
			c3                 => open,                                      --           (terminated)
			c4                 => open,                                      --           (terminated)
			areset             => '0',                                       --           (terminated)
			phasedone          => open,                                      --           (terminated)
			phasecounterselect => "000",                                     --           (terminated)
			phaseupdown        => '0',                                       --           (terminated)
			phasestep          => '0',                                       --           (terminated)
			scanclk            => '0',                                       --           (terminated)
			scanclkena         => '0',                                       --           (terminated)
			scandata           => '0',                                       --           (terminated)
			configupdate       => '0'                                        --           (terminated)
		);

	sdram_controller : component embedded_computer_system_sdram_controller
		port map (
			clk            => pll_c0_clk,                                                 --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,                   -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_controller_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_controller_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_controller_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_controller_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_controller_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_controller_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_controller_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_controller_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_controller_addr,                                      --  wire.export
			zs_ba          => sdram_controller_ba,                                        --      .export
			zs_cas_n       => sdram_controller_cas_n,                                     --      .export
			zs_cke         => sdram_controller_cke,                                       --      .export
			zs_cs_n        => sdram_controller_cs_n,                                      --      .export
			zs_dq          => sdram_controller_dq,                                        --      .export
			zs_dqm         => sdram_controller_dqm,                                       --      .export
			zs_ras_n       => sdram_controller_ras_n,                                     --      .export
			zs_we_n        => sdram_controller_we_n                                       --      .export
		);

	sierra_0 : component sierra
		port map (
			address                     => mm_interconnect_0_sierra_0_avalon_slave_0_address,              --    avalon_slave_0.address
			chipselect_n                => mm_interconnect_0_sierra_0_avalon_slave_0_chipselect_ports_inv, --                  .chipselect_n
			read_n                      => mm_interconnect_0_sierra_0_avalon_slave_0_read_ports_inv,       --                  .read_n
			writedata                   => mm_interconnect_0_sierra_0_avalon_slave_0_writedata,            --                  .writedata
			write_n                     => mm_interconnect_0_sierra_0_avalon_slave_0_write_ports_inv,      --                  .write_n
			readdata                    => mm_interconnect_0_sierra_0_avalon_slave_0_readdata,             --                  .readdata
			clk                         => pll_c0_clk,                                                     --       clock_reset.clk
			reset_n                     => rst_controller_001_reset_out_reset_ports_inv,                   -- clock_reset_reset.reset_n
			external_runing_taskid_info => sierra_0_conduit_end_export,                                    --       conduit_end.export
			irq                         => irq_mapper_receiver0_irq,                                       --  interrupt_sender.irq
			extirq_n                    => sierra_0_conduit_end_1_export                                   --     conduit_end_1.export
		);

	sysid_qsys_0 : component embedded_computer_system_sysid_qsys_0
		port map (
			clock    => pll_c0_clk,                                              --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	temperature_set_ip_0 : component temperature_set_IP
		port map (
			clk      => pll_c0_clk,                                                                 --          clock.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                                   --          reset.reset_n
			cs_n     => mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_chipselect_ports_inv, -- avalon_slave_0.chipselect_n
			read_n   => mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_read_ports_inv,       --               .read_n
			data_out => mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_readdata,             --               .readdata
			data_in  => temperature_set_ip_0_writedata                                              --    conduit_end.writedata
		);

	value_0 : component embedded_computer_system_value_0
		port map (
			avs_a_read         => mm_interconnect_0_value_0_avs_a_read,         --   avs_a.read
			avs_a_write        => mm_interconnect_0_value_0_avs_a_write,        --        .write
			avs_a_address      => mm_interconnect_0_value_0_avs_a_address,      --        .address
			avs_a_writedata    => mm_interconnect_0_value_0_avs_a_writedata,    --        .writedata
			avs_a_byteenable   => mm_interconnect_0_value_0_avs_a_byteenable,   --        .byteenable
			avs_a_readdata     => mm_interconnect_0_value_0_avs_a_readdata,     --        .readdata
			avs_cra_read       => mm_interconnect_0_value_0_avs_cra_read,       -- avs_cra.read
			avs_cra_write      => mm_interconnect_0_value_0_avs_cra_write,      --        .write
			avs_cra_address    => mm_interconnect_0_value_0_avs_cra_address,    --        .address
			avs_cra_writedata  => mm_interconnect_0_value_0_avs_cra_writedata,  --        .writedata
			avs_cra_byteenable => mm_interconnect_0_value_0_avs_cra_byteenable, --        .byteenable
			avs_cra_readdata   => mm_interconnect_0_value_0_avs_cra_readdata,   --        .readdata
			clock              => pll_c0_clk,                                   --   clock.clk
			done_irq           => irq_mapper_receiver2_irq,                     --     irq.irq
			resetn             => rst_controller_reset_out_reset_ports_inv      --   reset.reset_n
		);

	mm_interconnect_0 : component embedded_computer_system_mm_interconnect_0
		port map (
			clk_0_clk_clk                                         => clk_clk,                                                          --                                       clk_0_clk.clk
			pll_c0_clk                                            => pll_c0_clk,                                                       --                                          pll_c0.clk
			cpu_reset_reset_bridge_in_reset_reset                 => rst_controller_001_reset_out_reset,                               --                 cpu_reset_reset_bridge_in_reset.reset
			jtag_uart_reset_reset_bridge_in_reset_reset           => rst_controller_reset_out_reset,                                   --           jtag_uart_reset_reset_bridge_in_reset.reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_002_reset_out_reset,                               -- pll_inclk_interface_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                               => cpu_data_master_address,                                          --                                 cpu_data_master.address
			cpu_data_master_waitrequest                           => cpu_data_master_waitrequest,                                      --                                                .waitrequest
			cpu_data_master_byteenable                            => cpu_data_master_byteenable,                                       --                                                .byteenable
			cpu_data_master_read                                  => cpu_data_master_read,                                             --                                                .read
			cpu_data_master_readdata                              => cpu_data_master_readdata,                                         --                                                .readdata
			cpu_data_master_write                                 => cpu_data_master_write,                                            --                                                .write
			cpu_data_master_writedata                             => cpu_data_master_writedata,                                        --                                                .writedata
			cpu_data_master_debugaccess                           => cpu_data_master_debugaccess,                                      --                                                .debugaccess
			cpu_instruction_master_address                        => cpu_instruction_master_address,                                   --                          cpu_instruction_master.address
			cpu_instruction_master_waitrequest                    => cpu_instruction_master_waitrequest,                               --                                                .waitrequest
			cpu_instruction_master_read                           => cpu_instruction_master_read,                                      --                                                .read
			cpu_instruction_master_readdata                       => cpu_instruction_master_readdata,                                  --                                                .readdata
			cpu_debug_mem_slave_address                           => mm_interconnect_0_cpu_debug_mem_slave_address,                    --                             cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                             => mm_interconnect_0_cpu_debug_mem_slave_write,                      --                                                .write
			cpu_debug_mem_slave_read                              => mm_interconnect_0_cpu_debug_mem_slave_read,                       --                                                .read
			cpu_debug_mem_slave_readdata                          => mm_interconnect_0_cpu_debug_mem_slave_readdata,                   --                                                .readdata
			cpu_debug_mem_slave_writedata                         => mm_interconnect_0_cpu_debug_mem_slave_writedata,                  --                                                .writedata
			cpu_debug_mem_slave_byteenable                        => mm_interconnect_0_cpu_debug_mem_slave_byteenable,                 --                                                .byteenable
			cpu_debug_mem_slave_waitrequest                       => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,                --                                                .waitrequest
			cpu_debug_mem_slave_debugaccess                       => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,                --                                                .debugaccess
			jtag_uart_avalon_jtag_slave_address                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,            --                     jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,              --                                                .write
			jtag_uart_avalon_jtag_slave_read                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,               --                                                .read
			jtag_uart_avalon_jtag_slave_readdata                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,           --                                                .readdata
			jtag_uart_avalon_jtag_slave_writedata                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,          --                                                .writedata
			jtag_uart_avalon_jtag_slave_waitrequest               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,        --                                                .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,         --                                                .chipselect
			modular_adc_0_sample_store_csr_address                => mm_interconnect_0_modular_adc_0_sample_store_csr_address,         --                  modular_adc_0_sample_store_csr.address
			modular_adc_0_sample_store_csr_write                  => mm_interconnect_0_modular_adc_0_sample_store_csr_write,           --                                                .write
			modular_adc_0_sample_store_csr_read                   => mm_interconnect_0_modular_adc_0_sample_store_csr_read,            --                                                .read
			modular_adc_0_sample_store_csr_readdata               => mm_interconnect_0_modular_adc_0_sample_store_csr_readdata,        --                                                .readdata
			modular_adc_0_sample_store_csr_writedata              => mm_interconnect_0_modular_adc_0_sample_store_csr_writedata,       --                                                .writedata
			modular_adc_0_sequencer_csr_address                   => mm_interconnect_0_modular_adc_0_sequencer_csr_address,            --                     modular_adc_0_sequencer_csr.address
			modular_adc_0_sequencer_csr_write                     => mm_interconnect_0_modular_adc_0_sequencer_csr_write,              --                                                .write
			modular_adc_0_sequencer_csr_read                      => mm_interconnect_0_modular_adc_0_sequencer_csr_read,               --                                                .read
			modular_adc_0_sequencer_csr_readdata                  => mm_interconnect_0_modular_adc_0_sequencer_csr_readdata,           --                                                .readdata
			modular_adc_0_sequencer_csr_writedata                 => mm_interconnect_0_modular_adc_0_sequencer_csr_writedata,          --                                                .writedata
			pio_0_s1_address                                      => mm_interconnect_0_pio_0_s1_address,                               --                                        pio_0_s1.address
			pio_0_s1_write                                        => mm_interconnect_0_pio_0_s1_write,                                 --                                                .write
			pio_0_s1_readdata                                     => mm_interconnect_0_pio_0_s1_readdata,                              --                                                .readdata
			pio_0_s1_writedata                                    => mm_interconnect_0_pio_0_s1_writedata,                             --                                                .writedata
			pio_0_s1_chipselect                                   => mm_interconnect_0_pio_0_s1_chipselect,                            --                                                .chipselect
			pll_pll_slave_address                                 => mm_interconnect_0_pll_pll_slave_address,                          --                                   pll_pll_slave.address
			pll_pll_slave_write                                   => mm_interconnect_0_pll_pll_slave_write,                            --                                                .write
			pll_pll_slave_read                                    => mm_interconnect_0_pll_pll_slave_read,                             --                                                .read
			pll_pll_slave_readdata                                => mm_interconnect_0_pll_pll_slave_readdata,                         --                                                .readdata
			pll_pll_slave_writedata                               => mm_interconnect_0_pll_pll_slave_writedata,                        --                                                .writedata
			sdram_controller_s1_address                           => mm_interconnect_0_sdram_controller_s1_address,                    --                             sdram_controller_s1.address
			sdram_controller_s1_write                             => mm_interconnect_0_sdram_controller_s1_write,                      --                                                .write
			sdram_controller_s1_read                              => mm_interconnect_0_sdram_controller_s1_read,                       --                                                .read
			sdram_controller_s1_readdata                          => mm_interconnect_0_sdram_controller_s1_readdata,                   --                                                .readdata
			sdram_controller_s1_writedata                         => mm_interconnect_0_sdram_controller_s1_writedata,                  --                                                .writedata
			sdram_controller_s1_byteenable                        => mm_interconnect_0_sdram_controller_s1_byteenable,                 --                                                .byteenable
			sdram_controller_s1_readdatavalid                     => mm_interconnect_0_sdram_controller_s1_readdatavalid,              --                                                .readdatavalid
			sdram_controller_s1_waitrequest                       => mm_interconnect_0_sdram_controller_s1_waitrequest,                --                                                .waitrequest
			sdram_controller_s1_chipselect                        => mm_interconnect_0_sdram_controller_s1_chipselect,                 --                                                .chipselect
			sierra_0_avalon_slave_0_address                       => mm_interconnect_0_sierra_0_avalon_slave_0_address,                --                         sierra_0_avalon_slave_0.address
			sierra_0_avalon_slave_0_write                         => mm_interconnect_0_sierra_0_avalon_slave_0_write,                  --                                                .write
			sierra_0_avalon_slave_0_read                          => mm_interconnect_0_sierra_0_avalon_slave_0_read,                   --                                                .read
			sierra_0_avalon_slave_0_readdata                      => mm_interconnect_0_sierra_0_avalon_slave_0_readdata,               --                                                .readdata
			sierra_0_avalon_slave_0_writedata                     => mm_interconnect_0_sierra_0_avalon_slave_0_writedata,              --                                                .writedata
			sierra_0_avalon_slave_0_chipselect                    => mm_interconnect_0_sierra_0_avalon_slave_0_chipselect,             --                                                .chipselect
			sysid_qsys_0_control_slave_address                    => mm_interconnect_0_sysid_qsys_0_control_slave_address,             --                      sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                   => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,            --                                                .readdata
			temperature_set_IP_0_avalon_slave_0_read              => mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_read,       --             temperature_set_IP_0_avalon_slave_0.read
			temperature_set_IP_0_avalon_slave_0_readdata          => mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_readdata,   --                                                .readdata
			temperature_set_IP_0_avalon_slave_0_chipselect        => mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_chipselect, --                                                .chipselect
			value_0_avs_a_address                                 => mm_interconnect_0_value_0_avs_a_address,                          --                                   value_0_avs_a.address
			value_0_avs_a_write                                   => mm_interconnect_0_value_0_avs_a_write,                            --                                                .write
			value_0_avs_a_read                                    => mm_interconnect_0_value_0_avs_a_read,                             --                                                .read
			value_0_avs_a_readdata                                => mm_interconnect_0_value_0_avs_a_readdata,                         --                                                .readdata
			value_0_avs_a_writedata                               => mm_interconnect_0_value_0_avs_a_writedata,                        --                                                .writedata
			value_0_avs_a_byteenable                              => mm_interconnect_0_value_0_avs_a_byteenable,                       --                                                .byteenable
			value_0_avs_cra_address                               => mm_interconnect_0_value_0_avs_cra_address,                        --                                 value_0_avs_cra.address
			value_0_avs_cra_write                                 => mm_interconnect_0_value_0_avs_cra_write,                          --                                                .write
			value_0_avs_cra_read                                  => mm_interconnect_0_value_0_avs_cra_read,                           --                                                .read
			value_0_avs_cra_readdata                              => mm_interconnect_0_value_0_avs_cra_readdata,                       --                                                .readdata
			value_0_avs_cra_writedata                             => mm_interconnect_0_value_0_avs_cra_writedata,                      --                                                .writedata
			value_0_avs_cra_byteenable                            => mm_interconnect_0_value_0_avs_cra_byteenable,                     --                                                .byteenable
			VGA_IP_0_avalon_slave_0_address                       => mm_interconnect_0_vga_ip_0_avalon_slave_0_address,                --                         VGA_IP_0_avalon_slave_0.address
			VGA_IP_0_avalon_slave_0_write                         => mm_interconnect_0_vga_ip_0_avalon_slave_0_write,                  --                                                .write
			VGA_IP_0_avalon_slave_0_writedata                     => mm_interconnect_0_vga_ip_0_avalon_slave_0_writedata,              --                                                .writedata
			VGA_IP_0_avalon_slave_0_chipselect                    => mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect              --                                                .chipselect
		);

	irq_mapper : component embedded_computer_system_irq_mapper
		port map (
			clk           => pll_c0_clk,                         --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			sender_irq    => cpu_irq_irq                         --    sender.irq
		);

	rst_controller : component embedded_computer_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,        -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,  -- reset_in1.reset
			clk            => pll_c0_clk,                     --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component embedded_computer_system_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			clk            => pll_c0_clk,                             --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_in1      => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component embedded_computer_system_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect_ports_inv <= not mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect;

	mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_chipselect_ports_inv <= not mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_chipselect;

	mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_read_ports_inv <= not mm_interconnect_0_temperature_set_ip_0_avalon_slave_0_read;

	mm_interconnect_0_sierra_0_avalon_slave_0_chipselect_ports_inv <= not mm_interconnect_0_sierra_0_avalon_slave_0_chipselect;

	mm_interconnect_0_sierra_0_avalon_slave_0_read_ports_inv <= not mm_interconnect_0_sierra_0_avalon_slave_0_read;

	mm_interconnect_0_sierra_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_sierra_0_avalon_slave_0_write;

	mm_interconnect_0_sdram_controller_s1_read_ports_inv <= not mm_interconnect_0_sdram_controller_s1_read;

	mm_interconnect_0_sdram_controller_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_controller_s1_byteenable;

	mm_interconnect_0_sdram_controller_s1_write_ports_inv <= not mm_interconnect_0_sdram_controller_s1_write;

	mm_interconnect_0_pio_0_s1_write_ports_inv <= not mm_interconnect_0_pio_0_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of embedded_computer_system
