// tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module tb (
	);

	wire         clock_reset_inst_clock_clk;                                                                      // clock_reset_inst:clock -> [average_value_inst:clock, component_dpi_controller_average_value_inst:clock, irq_mapper:clk, main_dpi_controller_inst:clock, mm_interconnect_0:clock_reset_inst_clock_clk, mm_interconnect_1:clock_reset_inst_clock_clk, mm_master_dpi_bfm_average_value_avs_a_inst:clock, mm_master_dpi_bfm_average_value_avs_cra_inst:clock]
	wire         clock_reset_inst_clock2x_clk;                                                                    // clock_reset_inst:clock2x -> [component_dpi_controller_average_value_inst:clock2x, main_dpi_controller_inst:clock2x]
	wire         component_dpi_controller_average_value_inst_component_done_conduit;                              // component_dpi_controller_average_value_inst:component_done -> concatenate_component_done_inst:in_conduit_0
	wire   [0:0] main_dpi_controller_inst_component_enabled_conduit;                                              // main_dpi_controller_inst:component_enabled -> split_component_start_inst:in_conduit
	wire         component_dpi_controller_average_value_inst_component_wait_for_stream_writes_conduit;            // component_dpi_controller_average_value_inst:component_wait_for_stream_writes -> concatenate_component_wait_for_stream_writes_inst:in_conduit_0
	wire         mm_master_dpi_bfm_average_value_avs_a_inst_cra_control_done_writes_to_cra_conduit;               // mm_master_dpi_bfm_average_value_avs_a_inst:done_writes_to_cra -> average_value_component_cra_slave_memories_done_concatenate_inst:in_conduit_0
	wire         component_dpi_controller_average_value_inst_dpi_control_bind_conduit;                            // component_dpi_controller_average_value_inst:bind_interfaces -> average_value_component_dpi_controller_bind_conduit_fanout_inst:in_conduit
	wire         mm_master_dpi_bfm_average_value_avs_a_inst_dpi_control_done_reads_conduit;                       // mm_master_dpi_bfm_average_value_avs_a_inst:done_reads -> average_value_component_dpi_controller_slave_done_concatenate_inst:in_conduit_0
	wire         mm_master_dpi_bfm_average_value_avs_cra_inst_dpi_control_done_reads_conduit;                     // mm_master_dpi_bfm_average_value_avs_cra_inst:done_reads -> average_value_component_dpi_controller_slave_done_concatenate_inst:in_conduit_1
	wire         mm_master_dpi_bfm_average_value_avs_a_inst_dpi_control_done_writes_conduit;                      // mm_master_dpi_bfm_average_value_avs_a_inst:done_writes -> average_value_component_dpi_controller_slave_ready_concatenate_inst:in_conduit_0
	wire         mm_master_dpi_bfm_average_value_avs_cra_inst_dpi_control_done_writes_conduit;                    // mm_master_dpi_bfm_average_value_avs_cra_inst:done_writes -> average_value_component_dpi_controller_slave_ready_concatenate_inst:in_conduit_1
	wire         component_dpi_controller_average_value_inst_dpi_control_enable_conduit;                          // component_dpi_controller_average_value_inst:enable_interfaces -> average_value_component_dpi_controller_enable_conduit_fanout_inst:in_conduit
	wire         concatenate_component_done_inst_out_conduit_conduit;                                             // concatenate_component_done_inst:out_conduit -> main_dpi_controller_inst:component_done
	wire         concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit;                           // concatenate_component_wait_for_stream_writes_inst:out_conduit -> main_dpi_controller_inst:component_wait_for_stream_writes
	wire         average_value_component_cra_slave_memories_done_concatenate_inst_out_conduit_conduit;            // average_value_component_cra_slave_memories_done_concatenate_inst:out_conduit -> mm_master_dpi_bfm_average_value_avs_cra_inst:slave_memory_writes_done
	wire   [1:0] average_value_component_dpi_controller_slave_done_concatenate_inst_out_conduit_conduit;          // average_value_component_dpi_controller_slave_done_concatenate_inst:out_conduit -> component_dpi_controller_average_value_inst:slaves_done
	wire   [1:0] average_value_component_dpi_controller_slave_ready_concatenate_inst_out_conduit_conduit;         // average_value_component_dpi_controller_slave_ready_concatenate_inst:out_conduit -> component_dpi_controller_average_value_inst:slaves_ready
	wire         split_component_start_inst_out_conduit_0_conduit;                                                // split_component_start_inst:out_conduit_0 -> component_dpi_controller_average_value_inst:component_enabled
	wire         average_value_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit;           // average_value_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_0 -> mm_master_dpi_bfm_average_value_avs_a_inst:do_bind
	wire         average_value_component_dpi_controller_slave_readback_fanout_inst_out_conduit_0_conduit;         // average_value_component_dpi_controller_slave_readback_fanout_inst:out_conduit_0 -> mm_master_dpi_bfm_average_value_avs_a_inst:component_done
	wire         average_value_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit; // average_value_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_0 -> mm_master_dpi_bfm_average_value_avs_a_inst:component_started
	wire         average_value_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit;         // average_value_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_0 -> mm_master_dpi_bfm_average_value_avs_a_inst:enable
	wire         average_value_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit;           // average_value_component_dpi_controller_bind_conduit_fanout_inst:out_conduit_1 -> mm_master_dpi_bfm_average_value_avs_cra_inst:do_bind
	wire         average_value_component_dpi_controller_slave_readback_fanout_inst_out_conduit_1_conduit;         // average_value_component_dpi_controller_slave_readback_fanout_inst:out_conduit_1 -> mm_master_dpi_bfm_average_value_avs_cra_inst:component_done
	wire         average_value_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit; // average_value_component_dpi_controller_implicit_ready_conduit_fanout_inst:out_conduit_1 -> mm_master_dpi_bfm_average_value_avs_cra_inst:component_started
	wire         average_value_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit;         // average_value_component_dpi_controller_enable_conduit_fanout_inst:out_conduit_1 -> mm_master_dpi_bfm_average_value_avs_cra_inst:enable
	wire         component_dpi_controller_average_value_inst_read_implicit_streams_conduit;                       // component_dpi_controller_average_value_inst:read_implicit_streams -> average_value_component_dpi_controller_implicit_ready_conduit_fanout_inst:in_conduit
	wire         component_dpi_controller_average_value_inst_readback_from_slaves_conduit;                        // component_dpi_controller_average_value_inst:readback_from_slaves -> average_value_component_dpi_controller_slave_readback_fanout_inst:in_conduit
	wire         main_dpi_controller_inst_reset_ctrl_conduit;                                                     // main_dpi_controller_inst:trigger_reset -> clock_reset_inst:trigger_reset
	wire         clock_reset_inst_reset_reset;                                                                    // clock_reset_inst:resetn -> [average_value_inst:resetn, component_dpi_controller_average_value_inst:resetn, irq_mapper:reset, main_dpi_controller_inst:resetn, mm_interconnect_0:mm_master_dpi_bfm_average_value_avs_a_inst_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mm_master_dpi_bfm_average_value_avs_cra_inst_reset_reset_bridge_in_reset_reset, mm_master_dpi_bfm_average_value_avs_a_inst:reset_n, mm_master_dpi_bfm_average_value_avs_cra_inst:reset_n]
	wire   [7:0] mm_master_dpi_bfm_average_value_avs_a_inst_m0_readdata;                                          // mm_interconnect_0:mm_master_dpi_bfm_average_value_avs_a_inst_m0_readdata -> mm_master_dpi_bfm_average_value_avs_a_inst:avm_readdata
	wire         mm_master_dpi_bfm_average_value_avs_a_inst_m0_waitrequest;                                       // mm_interconnect_0:mm_master_dpi_bfm_average_value_avs_a_inst_m0_waitrequest -> mm_master_dpi_bfm_average_value_avs_a_inst:avm_waitrequest
	wire   [7:0] mm_master_dpi_bfm_average_value_avs_a_inst_m0_address;                                           // mm_master_dpi_bfm_average_value_avs_a_inst:avm_address -> mm_interconnect_0:mm_master_dpi_bfm_average_value_avs_a_inst_m0_address
	wire         mm_master_dpi_bfm_average_value_avs_a_inst_m0_read;                                              // mm_master_dpi_bfm_average_value_avs_a_inst:avm_read -> mm_interconnect_0:mm_master_dpi_bfm_average_value_avs_a_inst_m0_read
	wire   [0:0] mm_master_dpi_bfm_average_value_avs_a_inst_m0_byteenable;                                        // mm_master_dpi_bfm_average_value_avs_a_inst:avm_byteenable -> mm_interconnect_0:mm_master_dpi_bfm_average_value_avs_a_inst_m0_byteenable
	wire         mm_master_dpi_bfm_average_value_avs_a_inst_m0_readdatavalid;                                     // mm_interconnect_0:mm_master_dpi_bfm_average_value_avs_a_inst_m0_readdatavalid -> mm_master_dpi_bfm_average_value_avs_a_inst:avm_readdatavalid
	wire   [7:0] mm_master_dpi_bfm_average_value_avs_a_inst_m0_writedata;                                         // mm_master_dpi_bfm_average_value_avs_a_inst:avm_writedata -> mm_interconnect_0:mm_master_dpi_bfm_average_value_avs_a_inst_m0_writedata
	wire         mm_master_dpi_bfm_average_value_avs_a_inst_m0_write;                                             // mm_master_dpi_bfm_average_value_avs_a_inst:avm_write -> mm_interconnect_0:mm_master_dpi_bfm_average_value_avs_a_inst_m0_write
	wire   [0:0] mm_master_dpi_bfm_average_value_avs_a_inst_m0_burstcount;                                        // mm_master_dpi_bfm_average_value_avs_a_inst:avm_burstcount -> mm_interconnect_0:mm_master_dpi_bfm_average_value_avs_a_inst_m0_burstcount
	wire  [31:0] mm_interconnect_0_average_value_inst_avs_a_readdata;                                             // average_value_inst:avs_a_readdata -> mm_interconnect_0:average_value_inst_avs_a_readdata
	wire   [5:0] mm_interconnect_0_average_value_inst_avs_a_address;                                              // mm_interconnect_0:average_value_inst_avs_a_address -> average_value_inst:avs_a_address
	wire         mm_interconnect_0_average_value_inst_avs_a_read;                                                 // mm_interconnect_0:average_value_inst_avs_a_read -> average_value_inst:avs_a_read
	wire   [3:0] mm_interconnect_0_average_value_inst_avs_a_byteenable;                                           // mm_interconnect_0:average_value_inst_avs_a_byteenable -> average_value_inst:avs_a_byteenable
	wire         mm_interconnect_0_average_value_inst_avs_a_write;                                                // mm_interconnect_0:average_value_inst_avs_a_write -> average_value_inst:avs_a_write
	wire  [31:0] mm_interconnect_0_average_value_inst_avs_a_writedata;                                            // mm_interconnect_0:average_value_inst_avs_a_writedata -> average_value_inst:avs_a_writedata
	wire  [63:0] mm_master_dpi_bfm_average_value_avs_cra_inst_m0_readdata;                                        // mm_interconnect_1:mm_master_dpi_bfm_average_value_avs_cra_inst_m0_readdata -> mm_master_dpi_bfm_average_value_avs_cra_inst:avm_readdata
	wire         mm_master_dpi_bfm_average_value_avs_cra_inst_m0_waitrequest;                                     // mm_interconnect_1:mm_master_dpi_bfm_average_value_avs_cra_inst_m0_waitrequest -> mm_master_dpi_bfm_average_value_avs_cra_inst:avm_waitrequest
	wire   [5:0] mm_master_dpi_bfm_average_value_avs_cra_inst_m0_address;                                         // mm_master_dpi_bfm_average_value_avs_cra_inst:avm_address -> mm_interconnect_1:mm_master_dpi_bfm_average_value_avs_cra_inst_m0_address
	wire         mm_master_dpi_bfm_average_value_avs_cra_inst_m0_read;                                            // mm_master_dpi_bfm_average_value_avs_cra_inst:avm_read -> mm_interconnect_1:mm_master_dpi_bfm_average_value_avs_cra_inst_m0_read
	wire   [7:0] mm_master_dpi_bfm_average_value_avs_cra_inst_m0_byteenable;                                      // mm_master_dpi_bfm_average_value_avs_cra_inst:avm_byteenable -> mm_interconnect_1:mm_master_dpi_bfm_average_value_avs_cra_inst_m0_byteenable
	wire         mm_master_dpi_bfm_average_value_avs_cra_inst_m0_readdatavalid;                                   // mm_interconnect_1:mm_master_dpi_bfm_average_value_avs_cra_inst_m0_readdatavalid -> mm_master_dpi_bfm_average_value_avs_cra_inst:avm_readdatavalid
	wire  [63:0] mm_master_dpi_bfm_average_value_avs_cra_inst_m0_writedata;                                       // mm_master_dpi_bfm_average_value_avs_cra_inst:avm_writedata -> mm_interconnect_1:mm_master_dpi_bfm_average_value_avs_cra_inst_m0_writedata
	wire         mm_master_dpi_bfm_average_value_avs_cra_inst_m0_write;                                           // mm_master_dpi_bfm_average_value_avs_cra_inst:avm_write -> mm_interconnect_1:mm_master_dpi_bfm_average_value_avs_cra_inst_m0_write
	wire   [0:0] mm_master_dpi_bfm_average_value_avs_cra_inst_m0_burstcount;                                      // mm_master_dpi_bfm_average_value_avs_cra_inst:avm_burstcount -> mm_interconnect_1:mm_master_dpi_bfm_average_value_avs_cra_inst_m0_burstcount
	wire  [63:0] mm_interconnect_1_average_value_inst_avs_cra_readdata;                                           // average_value_inst:avs_cra_readdata -> mm_interconnect_1:average_value_inst_avs_cra_readdata
	wire   [2:0] mm_interconnect_1_average_value_inst_avs_cra_address;                                            // mm_interconnect_1:average_value_inst_avs_cra_address -> average_value_inst:avs_cra_address
	wire         mm_interconnect_1_average_value_inst_avs_cra_read;                                               // mm_interconnect_1:average_value_inst_avs_cra_read -> average_value_inst:avs_cra_read
	wire   [7:0] mm_interconnect_1_average_value_inst_avs_cra_byteenable;                                         // mm_interconnect_1:average_value_inst_avs_cra_byteenable -> average_value_inst:avs_cra_byteenable
	wire         mm_interconnect_1_average_value_inst_avs_cra_write;                                              // mm_interconnect_1:average_value_inst_avs_cra_write -> average_value_inst:avs_cra_write
	wire  [63:0] mm_interconnect_1_average_value_inst_avs_cra_writedata;                                          // mm_interconnect_1:average_value_inst_avs_cra_writedata -> average_value_inst:avs_cra_writedata
	wire         irq_mapper_receiver0_irq;                                                                        // average_value_inst:done_irq -> irq_mapper:receiver0_irq
	wire         component_dpi_controller_average_value_inst_component_irq_irq;                                   // irq_mapper:sender_irq -> component_dpi_controller_average_value_inst:done_irq

	tb_average_value_component_cra_slave_memories_done_concatenate_inst average_value_component_cra_slave_memories_done_concatenate_inst (
		.out_conduit  (average_value_component_cra_slave_memories_done_concatenate_inst_out_conduit_conduit), //  out_conduit.conduit
		.in_conduit_0 (mm_master_dpi_bfm_average_value_avs_a_inst_cra_control_done_writes_to_cra_conduit)     // in_conduit_0.conduit
	);

	tb_average_value_component_dpi_controller_bind_conduit_fanout_inst average_value_component_dpi_controller_bind_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_average_value_inst_dpi_control_bind_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (average_value_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (average_value_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit)  // out_conduit_1.conduit
	);

	tb_average_value_component_dpi_controller_bind_conduit_fanout_inst average_value_component_dpi_controller_enable_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_average_value_inst_dpi_control_enable_conduit),                  //    in_conduit.conduit
		.out_conduit_0 (average_value_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (average_value_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit)  // out_conduit_1.conduit
	);

	tb_average_value_component_dpi_controller_bind_conduit_fanout_inst average_value_component_dpi_controller_implicit_ready_conduit_fanout_inst (
		.in_conduit    (component_dpi_controller_average_value_inst_read_implicit_streams_conduit),                       //    in_conduit.conduit
		.out_conduit_0 (average_value_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (average_value_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit)  // out_conduit_1.conduit
	);

	tb_average_value_component_dpi_controller_slave_done_concatenate_inst average_value_component_dpi_controller_slave_done_concatenate_inst (
		.out_conduit  (average_value_component_dpi_controller_slave_done_concatenate_inst_out_conduit_conduit), //  out_conduit.conduit
		.in_conduit_0 (mm_master_dpi_bfm_average_value_avs_a_inst_dpi_control_done_reads_conduit),              // in_conduit_0.conduit
		.in_conduit_1 (mm_master_dpi_bfm_average_value_avs_cra_inst_dpi_control_done_reads_conduit)             // in_conduit_1.conduit
	);

	tb_average_value_component_dpi_controller_bind_conduit_fanout_inst average_value_component_dpi_controller_slave_readback_fanout_inst (
		.in_conduit    (component_dpi_controller_average_value_inst_readback_from_slaves_conduit),                //    in_conduit.conduit
		.out_conduit_0 (average_value_component_dpi_controller_slave_readback_fanout_inst_out_conduit_0_conduit), // out_conduit_0.conduit
		.out_conduit_1 (average_value_component_dpi_controller_slave_readback_fanout_inst_out_conduit_1_conduit)  // out_conduit_1.conduit
	);

	tb_average_value_component_dpi_controller_slave_done_concatenate_inst average_value_component_dpi_controller_slave_ready_concatenate_inst (
		.out_conduit  (average_value_component_dpi_controller_slave_ready_concatenate_inst_out_conduit_conduit), //  out_conduit.conduit
		.in_conduit_0 (mm_master_dpi_bfm_average_value_avs_a_inst_dpi_control_done_writes_conduit),              // in_conduit_0.conduit
		.in_conduit_1 (mm_master_dpi_bfm_average_value_avs_cra_inst_dpi_control_done_writes_conduit)             // in_conduit_1.conduit
	);

	tb_average_value_inst average_value_inst (
		.avs_a_read         (mm_interconnect_0_average_value_inst_avs_a_read),         //   avs_a.read
		.avs_a_write        (mm_interconnect_0_average_value_inst_avs_a_write),        //        .write
		.avs_a_address      (mm_interconnect_0_average_value_inst_avs_a_address),      //        .address
		.avs_a_writedata    (mm_interconnect_0_average_value_inst_avs_a_writedata),    //        .writedata
		.avs_a_byteenable   (mm_interconnect_0_average_value_inst_avs_a_byteenable),   //        .byteenable
		.avs_a_readdata     (mm_interconnect_0_average_value_inst_avs_a_readdata),     //        .readdata
		.avs_cra_read       (mm_interconnect_1_average_value_inst_avs_cra_read),       // avs_cra.read
		.avs_cra_write      (mm_interconnect_1_average_value_inst_avs_cra_write),      //        .write
		.avs_cra_address    (mm_interconnect_1_average_value_inst_avs_cra_address),    //        .address
		.avs_cra_writedata  (mm_interconnect_1_average_value_inst_avs_cra_writedata),  //        .writedata
		.avs_cra_byteenable (mm_interconnect_1_average_value_inst_avs_cra_byteenable), //        .byteenable
		.avs_cra_readdata   (mm_interconnect_1_average_value_inst_avs_cra_readdata),   //        .readdata
		.clock              (clock_reset_inst_clock_clk),                              //   clock.clk
		.done_irq           (irq_mapper_receiver0_irq),                                //     irq.irq
		.resetn             (clock_reset_inst_reset_reset)                             //   reset.reset_n
	);

	hls_sim_clock_reset #(
		.RESET_CYCLE_HOLD (4)
	) clock_reset_inst (
		.clock         (clock_reset_inst_clock_clk),                  //      clock.clk
		.resetn        (clock_reset_inst_reset_reset),                //      reset.reset_n
		.clock2x       (clock_reset_inst_clock2x_clk),                //    clock2x.clk
		.trigger_reset (main_dpi_controller_inst_reset_ctrl_conduit)  // reset_ctrl.conduit
	);

	hls_sim_component_dpi_controller #(
		.COMPONENT_NAME               ("average_value"),
		.RETURN_DATAWIDTH             (64),
		.COMPONENT_NUM_SLAVES         (2),
		.COMPONENT_HAS_SLAVE_RETURN   (1),
		.COMPONENT_NUM_OUTPUT_STREAMS (0)
	) component_dpi_controller_average_value_inst (
		.clock                            (clock_reset_inst_clock_clk),                                                              //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                                            //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                                            //                          clock2x.clk
		.bind_interfaces                  (component_dpi_controller_average_value_inst_dpi_control_bind_conduit),                    //                 dpi_control_bind.conduit
		.enable_interfaces                (component_dpi_controller_average_value_inst_dpi_control_enable_conduit),                  //               dpi_control_enable.conduit
		.slaves_ready                     (average_value_component_dpi_controller_slave_ready_concatenate_inst_out_conduit_conduit), //         dpi_control_slaves_ready.conduit
		.slaves_done                      (average_value_component_dpi_controller_slave_done_concatenate_inst_out_conduit_conduit),  //          dpi_control_slaves_done.conduit
		.component_enabled                (split_component_start_inst_out_conduit_0_conduit),                                        //                component_enabled.conduit
		.component_done                   (component_dpi_controller_average_value_inst_component_done_conduit),                      //                   component_done.conduit
		.component_wait_for_stream_writes (component_dpi_controller_average_value_inst_component_wait_for_stream_writes_conduit),    // component_wait_for_stream_writes.conduit
		.read_implicit_streams            (component_dpi_controller_average_value_inst_read_implicit_streams_conduit),               //            read_implicit_streams.conduit
		.readback_from_slaves             (component_dpi_controller_average_value_inst_readback_from_slaves_conduit),                //             readback_from_slaves.conduit
		.start                            (),                                                                                        //                   component_call.valid
		.done                             (),                                                                                        //                 component_return.valid
		.stall                            (),                                                                                        //                                 .stall
		.done_irq                         (component_dpi_controller_average_value_inst_component_irq_irq),                           //                    component_irq.irq
		.returndata                       (),                                                                                        //                       returndata.data
		.busy                             (1'b0)                                                                                     //                      (terminated)
	);

	tb_average_value_component_cra_slave_memories_done_concatenate_inst concatenate_component_done_inst (
		.out_conduit  (concatenate_component_done_inst_out_conduit_conduit),                //  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_average_value_inst_component_done_conduit)  // in_conduit_0.conduit
	);

	tb_average_value_component_cra_slave_memories_done_concatenate_inst concatenate_component_wait_for_stream_writes_inst (
		.out_conduit  (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit),                //  out_conduit.conduit
		.in_conduit_0 (component_dpi_controller_average_value_inst_component_wait_for_stream_writes_conduit)  // in_conduit_0.conduit
	);

	hls_sim_main_dpi_controller #(
		.NUM_COMPONENTS      (1),
		.COMPONENT_NAMES_STR ("average_value")
	) main_dpi_controller_inst (
		.clock                            (clock_reset_inst_clock_clk),                                            //                            clock.clk
		.resetn                           (clock_reset_inst_reset_reset),                                          //                            reset.reset_n
		.clock2x                          (clock_reset_inst_clock2x_clk),                                          //                          clock2x.clk
		.component_enabled                (main_dpi_controller_inst_component_enabled_conduit),                    //                component_enabled.conduit
		.component_done                   (concatenate_component_done_inst_out_conduit_conduit),                   //                   component_done.conduit
		.component_wait_for_stream_writes (concatenate_component_wait_for_stream_writes_inst_out_conduit_conduit), // component_wait_for_stream_writes.conduit
		.trigger_reset                    (main_dpi_controller_inst_reset_ctrl_conduit)                            //                       reset_ctrl.conduit
	);

	hls_sim_mm_master_dpi_bfm #(
		.AV_ADDRESS_W                         (8),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (1),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (3),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("average_value"),
		.COMPONENT_HAS_SLAVE_RETURN           (0),
		.COMPONENT_SLAVE_WRITE_INTERFACE_NAME ("a"),
		.COMPONENT_SLAVE_READ_INTERFACE_NAME  ("a_avs_readback"),
		.COMPONENT_CRA_SLAVE                  (0),
		.NUM_SLAVE_MEMORIES                   (0)
	) mm_master_dpi_bfm_average_value_avs_a_inst (
		.clock              (clock_reset_inst_clock_clk),                                                                      //                          clock.clk
		.reset_n            (clock_reset_inst_reset_reset),                                                                    //                          reset.reset_n
		.do_bind            (average_value_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_0_conduit),           //               dpi_control_bind.conduit
		.enable             (average_value_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_0_conduit),         //             dpi_control_enable.conduit
		.done_writes        (mm_master_dpi_bfm_average_value_avs_a_inst_dpi_control_done_writes_conduit),                      //        dpi_control_done_writes.conduit
		.done_reads         (mm_master_dpi_bfm_average_value_avs_a_inst_dpi_control_done_reads_conduit),                       //         dpi_control_done_reads.conduit
		.component_started  (average_value_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_0_conduit), //  dpi_control_component_started.conduit
		.component_done     (average_value_component_dpi_controller_slave_readback_fanout_inst_out_conduit_0_conduit),         //     dpi_control_component_done.conduit
		.done_writes_to_cra (mm_master_dpi_bfm_average_value_avs_a_inst_cra_control_done_writes_to_cra_conduit),               // cra_control_done_writes_to_cra.conduit
		.avm_writedata      (mm_master_dpi_bfm_average_value_avs_a_inst_m0_writedata),                                         //                             m0.writedata
		.avm_burstcount     (mm_master_dpi_bfm_average_value_avs_a_inst_m0_burstcount),                                        //                               .burstcount
		.avm_readdata       (mm_master_dpi_bfm_average_value_avs_a_inst_m0_readdata),                                          //                               .readdata
		.avm_address        (mm_master_dpi_bfm_average_value_avs_a_inst_m0_address),                                           //                               .address
		.avm_waitrequest    (mm_master_dpi_bfm_average_value_avs_a_inst_m0_waitrequest),                                       //                               .waitrequest
		.avm_write          (mm_master_dpi_bfm_average_value_avs_a_inst_m0_write),                                             //                               .write
		.avm_read           (mm_master_dpi_bfm_average_value_avs_a_inst_m0_read),                                              //                               .read
		.avm_byteenable     (mm_master_dpi_bfm_average_value_avs_a_inst_m0_byteenable),                                        //                               .byteenable
		.avm_readdatavalid  (mm_master_dpi_bfm_average_value_avs_a_inst_m0_readdatavalid)                                      //                               .readdatavalid
	);

	hls_sim_mm_master_dpi_bfm #(
		.AV_ADDRESS_W                         (6),
		.AV_SYMBOL_W                          (8),
		.AV_NUMSYMBOLS                        (8),
		.AV_BURSTCOUNT_W                      (1),
		.USE_READ                             (1),
		.USE_WRITE                            (1),
		.USE_ADDRESS                          (1),
		.USE_BYTE_ENABLE                      (1),
		.USE_BURSTCOUNT                       (0),
		.USE_READ_DATA                        (1),
		.USE_READ_DATA_VALID                  (1),
		.USE_WRITE_DATA                       (1),
		.USE_BEGIN_TRANSFER                   (0),
		.USE_BEGIN_BURST_TRANSFER             (0),
		.USE_WAIT_REQUEST                     (1),
		.AV_BURST_LINEWRAP                    (1),
		.AV_BURST_BNDR_ONLY                   (1),
		.AV_FIX_READ_LATENCY                  (1),
		.AV_READ_WAIT_TIME                    (0),
		.AV_WRITE_WAIT_TIME                   (0),
		.REGISTER_WAITREQUEST                 (0),
		.AV_REGISTERINCOMINGSIGNALS           (0),
		.COMPONENT_NAME                       ("average_value"),
		.COMPONENT_HAS_SLAVE_RETURN           (1),
		.COMPONENT_SLAVE_WRITE_INTERFACE_NAME ("__ihc_hls_avs_write_stream__"),
		.COMPONENT_SLAVE_READ_INTERFACE_NAME  ("$return"),
		.COMPONENT_CRA_SLAVE                  (1),
		.NUM_SLAVE_MEMORIES                   (1)
	) mm_master_dpi_bfm_average_value_avs_cra_inst (
		.clock                    (clock_reset_inst_clock_clk),                                                                      //                                clock.clk
		.reset_n                  (clock_reset_inst_reset_reset),                                                                    //                                reset.reset_n
		.do_bind                  (average_value_component_dpi_controller_bind_conduit_fanout_inst_out_conduit_1_conduit),           //                     dpi_control_bind.conduit
		.enable                   (average_value_component_dpi_controller_enable_conduit_fanout_inst_out_conduit_1_conduit),         //                   dpi_control_enable.conduit
		.done_writes              (mm_master_dpi_bfm_average_value_avs_cra_inst_dpi_control_done_writes_conduit),                    //              dpi_control_done_writes.conduit
		.done_reads               (mm_master_dpi_bfm_average_value_avs_cra_inst_dpi_control_done_reads_conduit),                     //               dpi_control_done_reads.conduit
		.component_started        (average_value_component_dpi_controller_implicit_ready_conduit_fanout_inst_out_conduit_1_conduit), //        dpi_control_component_started.conduit
		.component_done           (average_value_component_dpi_controller_slave_readback_fanout_inst_out_conduit_1_conduit),         //           dpi_control_component_done.conduit
		.done_writes_to_cra       (),                                                                                                //       cra_control_done_writes_to_cra.conduit
		.slave_memory_writes_done (average_value_component_cra_slave_memories_done_concatenate_inst_out_conduit_conduit),            // cra_control_slave_memory_writes_done.conduit
		.avm_writedata            (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_writedata),                                       //                                   m0.writedata
		.avm_burstcount           (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_burstcount),                                      //                                     .burstcount
		.avm_readdata             (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_readdata),                                        //                                     .readdata
		.avm_address              (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_address),                                         //                                     .address
		.avm_waitrequest          (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_waitrequest),                                     //                                     .waitrequest
		.avm_write                (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_write),                                           //                                     .write
		.avm_read                 (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_read),                                            //                                     .read
		.avm_byteenable           (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_byteenable),                                      //                                     .byteenable
		.avm_readdatavalid        (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_readdatavalid)                                    //                                     .readdatavalid
	);

	tb_split_component_start_inst split_component_start_inst (
		.in_conduit    (main_dpi_controller_inst_component_enabled_conduit), //    in_conduit.conduit
		.out_conduit_0 (split_component_start_inst_out_conduit_0_conduit)    // out_conduit_0.conduit
	);

	tb_mm_interconnect_0 mm_interconnect_0 (
		.clock_reset_inst_clock_clk                                                   (clock_reset_inst_clock_clk),                                  //                                                 clock_reset_inst_clock.clk
		.mm_master_dpi_bfm_average_value_avs_a_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                               // mm_master_dpi_bfm_average_value_avs_a_inst_reset_reset_bridge_in_reset.reset
		.mm_master_dpi_bfm_average_value_avs_a_inst_m0_address                        (mm_master_dpi_bfm_average_value_avs_a_inst_m0_address),       //                          mm_master_dpi_bfm_average_value_avs_a_inst_m0.address
		.mm_master_dpi_bfm_average_value_avs_a_inst_m0_waitrequest                    (mm_master_dpi_bfm_average_value_avs_a_inst_m0_waitrequest),   //                                                                       .waitrequest
		.mm_master_dpi_bfm_average_value_avs_a_inst_m0_burstcount                     (mm_master_dpi_bfm_average_value_avs_a_inst_m0_burstcount),    //                                                                       .burstcount
		.mm_master_dpi_bfm_average_value_avs_a_inst_m0_byteenable                     (mm_master_dpi_bfm_average_value_avs_a_inst_m0_byteenable),    //                                                                       .byteenable
		.mm_master_dpi_bfm_average_value_avs_a_inst_m0_read                           (mm_master_dpi_bfm_average_value_avs_a_inst_m0_read),          //                                                                       .read
		.mm_master_dpi_bfm_average_value_avs_a_inst_m0_readdata                       (mm_master_dpi_bfm_average_value_avs_a_inst_m0_readdata),      //                                                                       .readdata
		.mm_master_dpi_bfm_average_value_avs_a_inst_m0_readdatavalid                  (mm_master_dpi_bfm_average_value_avs_a_inst_m0_readdatavalid), //                                                                       .readdatavalid
		.mm_master_dpi_bfm_average_value_avs_a_inst_m0_write                          (mm_master_dpi_bfm_average_value_avs_a_inst_m0_write),         //                                                                       .write
		.mm_master_dpi_bfm_average_value_avs_a_inst_m0_writedata                      (mm_master_dpi_bfm_average_value_avs_a_inst_m0_writedata),     //                                                                       .writedata
		.average_value_inst_avs_a_address                                             (mm_interconnect_0_average_value_inst_avs_a_address),          //                                               average_value_inst_avs_a.address
		.average_value_inst_avs_a_write                                               (mm_interconnect_0_average_value_inst_avs_a_write),            //                                                                       .write
		.average_value_inst_avs_a_read                                                (mm_interconnect_0_average_value_inst_avs_a_read),             //                                                                       .read
		.average_value_inst_avs_a_readdata                                            (mm_interconnect_0_average_value_inst_avs_a_readdata),         //                                                                       .readdata
		.average_value_inst_avs_a_writedata                                           (mm_interconnect_0_average_value_inst_avs_a_writedata),        //                                                                       .writedata
		.average_value_inst_avs_a_byteenable                                          (mm_interconnect_0_average_value_inst_avs_a_byteenable)        //                                                                       .byteenable
	);

	tb_mm_interconnect_1 mm_interconnect_1 (
		.clock_reset_inst_clock_clk                                                     (clock_reset_inst_clock_clk),                                    //                                                   clock_reset_inst_clock.clk
		.mm_master_dpi_bfm_average_value_avs_cra_inst_reset_reset_bridge_in_reset_reset (~clock_reset_inst_reset_reset),                                 // mm_master_dpi_bfm_average_value_avs_cra_inst_reset_reset_bridge_in_reset.reset
		.mm_master_dpi_bfm_average_value_avs_cra_inst_m0_address                        (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_address),       //                          mm_master_dpi_bfm_average_value_avs_cra_inst_m0.address
		.mm_master_dpi_bfm_average_value_avs_cra_inst_m0_waitrequest                    (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_waitrequest),   //                                                                         .waitrequest
		.mm_master_dpi_bfm_average_value_avs_cra_inst_m0_burstcount                     (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_burstcount),    //                                                                         .burstcount
		.mm_master_dpi_bfm_average_value_avs_cra_inst_m0_byteenable                     (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_byteenable),    //                                                                         .byteenable
		.mm_master_dpi_bfm_average_value_avs_cra_inst_m0_read                           (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_read),          //                                                                         .read
		.mm_master_dpi_bfm_average_value_avs_cra_inst_m0_readdata                       (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_readdata),      //                                                                         .readdata
		.mm_master_dpi_bfm_average_value_avs_cra_inst_m0_readdatavalid                  (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_readdatavalid), //                                                                         .readdatavalid
		.mm_master_dpi_bfm_average_value_avs_cra_inst_m0_write                          (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_write),         //                                                                         .write
		.mm_master_dpi_bfm_average_value_avs_cra_inst_m0_writedata                      (mm_master_dpi_bfm_average_value_avs_cra_inst_m0_writedata),     //                                                                         .writedata
		.average_value_inst_avs_cra_address                                             (mm_interconnect_1_average_value_inst_avs_cra_address),          //                                               average_value_inst_avs_cra.address
		.average_value_inst_avs_cra_write                                               (mm_interconnect_1_average_value_inst_avs_cra_write),            //                                                                         .write
		.average_value_inst_avs_cra_read                                                (mm_interconnect_1_average_value_inst_avs_cra_read),             //                                                                         .read
		.average_value_inst_avs_cra_readdata                                            (mm_interconnect_1_average_value_inst_avs_cra_readdata),         //                                                                         .readdata
		.average_value_inst_avs_cra_writedata                                           (mm_interconnect_1_average_value_inst_avs_cra_writedata),        //                                                                         .writedata
		.average_value_inst_avs_cra_byteenable                                          (mm_interconnect_1_average_value_inst_avs_cra_byteenable)        //                                                                         .byteenable
	);

	tb_irq_mapper irq_mapper (
		.clk           (clock_reset_inst_clock_clk),                                    //       clk.clk
		.reset         (~clock_reset_inst_reset_reset),                                 // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),                                      // receiver0.irq
		.sender_irq    (component_dpi_controller_average_value_inst_component_irq_irq)  //    sender.irq
	);

endmodule
