��/  ���t\����h(u�;����u|q�ak�Ӷs�J������M��=�Ii�	T|}���\�pq��d|J"�n��1j�30��ڢ �@����)w�U�R�s�I��<;�
��\�xZ0�L�=g�Xl!`����L���u��X+}�ݰ��!^�0d��o߹���ɯyw:=G�`�9�PyCE��8%X�7	]�*����pogU��(~X� ��Vrv����P�Uh:l���V�	�$���p�2��_1y�ȯ�u� 4�D�M��hݿDI� 6�pn�l�!`' ��-1�=<H_6�n����(
'��UE��_Y2�&?�8dF��\��K�6� �y�滽4��b��[��d%����\Q�/�A�g�궷��Q��PTT�,/l[�fo+�)�2�~]牠�|��y�8���.c������� ���\���E�W��y[Y1Ԭ.��Μ�GSm?щn��K@F�R}q���#`/�?�㵵-+	��P�V��ñԷ"j(�]�Z��G4Ǌ���<�طX5��d�9�O%�F�9R6��1�w/�W?��^�K�7-�_b��0��X��7M����X��QH{G�Q�G���z���,z��ul5�Q7����G�o�؈�\���{j�NI���t;0��uE��w~�}0#g�ސ��I�y������|=:�B7���PHA���y0:�$a�{p�@��mB�(Ȓ��`�Ih�����G������7�)~DQ��2�46��eG2��7���������XL��&h���e���a_�cD������N7ٸ�c�m��j�����G�
嫙	Wxk#Oa�q
��e�b1]�$�<p��6�X�[��ئ���L�?�)t:��Y�/��U�O�Z�|E���]a��t��p���7Dk�r����ʬ�e���T��&��$���̡?;��t��-��y��yZ�Υ��}E�{���R�~��Nz����q,߄e	,�<��U]f�	��l|MO��q��n&SMb�^;�w{�s�7���@�LfBX�!H�XLQ^]��q����'eX�g�u�%�%e�f�'Q!�2�W���u�u3��wPm�������������}G�ג��<���+[��R?�ۊ&��*I�&�<�����>vjя�ȕ��Ԭ��ͺ��Z�>(�Ρ�T�ޒ�Ŗ�]�'�7�8�G��t0D⟽�����ݭ���1�_���ҡ�z7M�Ƅ{�%�]c��O̎P�):y|�e*��=9�>��X�uڅ�9�hՁ��������^!T��4@/I���z�(Q���:�����|ȁ�]T�V=�K��"��'&�+\�۪�N�G���L2���^Rq�����Fv\S�k�/`�R��
����=���fۈ��m>DN��!^s;^+�����J�@��V/�7���ycUSQ���:�R�v^9�'�kd�{/�Q�9<�����P���{�L#�h��a���,,'�{�k
���Xdr���j���V|�MT���磘�%j;Ğ����HN��b�H�m��6�d ��s��c�J�F�A$!�7����Ά��R��,��T2��X!XB^P��!s���5��{�n���J�\�t~�\��'��a��hg�[�gƘ뢇�S��ֲ`���~���(��f7�*��0}v���d�q
�R��O�q��p+8_>���S�O���6�"���qz�z�Ӄ݈��!TKi�aOm'�������]'h����i=i��d�>�=b�T:�ϙ�&v�ɛ�%��5 �{;k����%?�ES���<��f�@�FR�]8MR6�r�����e��3`l�'��7?��xۍ��.|V7ˣ�9��Ԡ�H���Q���0~��<(�<�2[�x�X&�v+C����3�4��=_���S�l���^d��U�hC��簐������鿟��Pǵ�{l�2���h��?�F���ʶ9���R��ǥA���c�8�z'~r�	�X}r\EB�p��+�w�;u�NR�]];z�"�O�&�)+SV�$�^_�ش��қ�% i��D��.���[/��p�J�O��z��]�����` %o��xN~�#� ۝���4��H���E�����CƏK9 6��e�Prf'_k�P/�����S~��-�w0���T����ay	��Wl.|����\��m5��e)���� �kTB�8˛�c
��j��.9"
�T��3����/�r<�fu�̐a[�dGU�	UaD�	͖2D�ض��ܭ�U�n�ʤ���aj#	����F�Q�$q�yX<I���ߠ�!� ��6i�B��i�i��t�dvV�F��M&MoJs��Y��I�Ev ^*��m�jU�ٛ���6�7�4o�3JN��
�d�4<�4��=��<��?�ӰFjh�e�B�<�!�dZ�J�C��T Rǔ&SY'��Uqj��]���vh5�������qs��8�#~A@������L��A�yug�kh��$C�]3�CE�B٤~��:hO�u��Q�2kC��UA���'��lB�(@�59P��ҀK7S����������`�nX��i�ǡ5S�4�96�����8ƞNp��Xpsܪ�����M�+9 �q�^顝A���o���dɞ~*UonE}}�p���-[:9�����k��?%M>�f��;x9v�F��ϓ��q��2�U�`H Pw�*�+4��`YR '�<Vd�f�2�����0�#�1+�+/R�[u�����
L
�h�> r�Ε�Y����Jn�ov��aE��9�.8��(ei݃>�V�e�0ڒ0an��E�LeǙ���xґȮ�NQ�S3i��h�?|��~`} lD�ג�����E��n��",Ԩ&,�.����$��d5Km�*u����n�&l�<�(ߐ]N^qTw�#re��8�iD�ꫨɅ���m�7�.A8>�G����᪭���d))�ބ�0��OPԲ���Hu�oQz��&GTn�Tk��O�r���@d�.ŐD-#��4���>�����x�R����0��	���o���#�rL���S�~ie�8�CHH�W����D#ˍvp��Y���aX��	�� U��x��?�o��A��P�{�
d�b�7�Q�X��I�,Gĸ�Z#[ �(^����^�}(ǯ��4��Z֕��+
�]Bx�T���w�F#xdJ^EC��� �gTW��)�1�܄$)��A3�����D���W
2�d��ŝ���"-��9��6>���FG>єz�.�6�͂��
�6d�����1�ǜ/�{t�bڰ,V��R9�`�r�񎣏���d�T��ӊ����V��6G.�Z�X��1i�Yx�Oݻ}l5w�h�o�|�R�>��_;,��r�������2���}�s~)�[�&���`)�Kͳ�|�V,@�}�&�&���v2���7�q�DX���i�cR(��b�Ϩ�ժ3�ïѹ3L.��h۳�+�������p&�H�	FqVh^�$dȋ�a�� ,��l���^�k����#��s5O�^�8��� y #$�}x���zʸGW��q����*ͱh�Uo�N�㐇��n�H&��FF�'R3ynw�L5g�=��5�VԂ]��6�/���<�J�D�2�µ8�ACj��F�� r\��$K,��;��?�]�0��F>�4�u�7H=c��|9�����U ]]�皱�{@�# �S�!�Jm���6j�E���aNRc���(9^��x�5ӻb/ �	�󍉪�'&pc��`�
��1����b���HT�7}��.�L�RJ]�nޚ�,ۭ�Qc��	Lp":=;<��7�Hi�b-��r��_R4#]�J7�"&�0��	g�ש�[��5���,�j�~��!�\���0���Mm�)h�wP+i��D%�\�=S�^�5It6�°�?�Mԓ���:#��\O�8��&��h%��'���n6x.���͉�K:h?if&W���H�R�!���9z��Ht��D�~&$�SЅ�IHg�[g��S�BU\��y<TM�����q��"�f��V����s�H��� �Z�[a�ך���1�!���Ǫ'���p�ׂeM�wN�.�5��	Q����`+
��0:��$���T/+��im�dž\��B8ȳ�jYU����-N��ç��#<ٸ�&|V��s}�V ~���&z��,�Zo��7�?u�[H�K�`���� t�G�!шD��f-^����\�f&�<"a/ ��7򰠊$d�N:�tA�o���2^���A����č�2��+=����(��%eO����OuѸ��J;�f(�@�̐�$g�y�yD�Z���w?���ɍ��r��j�Y@�K.�T_ڵ����U����F�&������	i�_4Y\�R=�@ߵ
��z�APT	�%�P�N3�C���SP���§B��S�9G"#����p�A�F�NEXP�\-&ocg1��/ۍ�@5��T�,��m��WT��ID�Y��DJ$���F���ͧ~r��|��� ��F1&�|�yTߺ�՞"���w��H/
lteW9��h7�ևڟ5� �
�Ly�I��k��=�t�V�ࠌ����oA��1���>Of{qƔ�.�������'��Q!̞����å�b�����Cw����xѮJ�tHŵ�r�,� F���.!����~@���0�^���Da��I�#D�]�nsÅ��{��޲+��;��CL��k�*>k��H��H}ȜH�����4��@�)H��)�P[��x��3	���<�Z��b�r�A���H�ZY>!¸�]'���/���Qs~�+����K��~�n��T��Tk^D"�W]CO];�u��Ҁ�`�O�?\םĆ�����w7J
� .8\��+z��UCjA��31��>�0Jc�D��,p�~E�9��Z��$,|
��m��xF��hU]�#&v�6�?`��3��iV�u���)�+���?�g�uD�8�6R�}�8$��'�eW�WZ�Lv;����+������s�����6��E�*W婬r�<Rc5������F�X�I3�.ti��*r4Z���i��"�
zϫZ�Z�|L2���cQ� �m^2����VJގ�apUMY�F:`c45P,[�XW3*q���W�U4 ��FçL1��m`�X�Ar����Zq'v�(���V��,U�E��0hҤ��G<4���*��C�Dш��ݙ��aGk�R1>��W�e��.��S5�Qj����'`~̂O<t�Xi-(�h��3�+�����1t2u��L;��ވ]́G�ϵ(̨s�z�D�d�,�f��^����4k���g�y_��S5�	e&I�f=�K�@�/��ܣ:���l�'oOs���;�����\���}l�я��B�|?7�	���&�sT����rK�X�p�P�Ks٘�[2��*E�y�=��˻��!�`������U������R�+��;��5���;��]Ý��Q�v���l����aGe����������$��cT��Qȸ�S���َ����Т�*����\����@>�WWc��A��#����X�.OQ��%rI�����d�n!� ��:���C;�we��5P��G%?��WY�.p	�f�C���P�^T_<�F���Ѯ�Œ���C!@���Ux7�0��1�qG����9�����?/y"�s%���[��c�;�п�s:^`L��aP�8ڔ�wQ��UN=�����d���U�C� -�vtĐ��f5ع�Id�k��D �b^��b� �D��.�y���oE�46h�֤��h��� Ƶ3:n.�A����'�eq��>ն�6�d5��?:|��â�����y[;C���c�h�ၥ
ӧcq@�Ν��SP\]˂���)�6!`|��h��⳷t�����\�c�����(nb�AE�����0�2Peh��v�>20X/E;"�>���m��}1M0�����h����x��.�n�U���'��S��? e����h�1�f�����Q8[������Wfr�9b��aq��'P*���UK���a�z��v�u�Z��Z�}G��mC�Ξ��+�����/6�;���x9"N'�����"d��f�ER���-9ۗ����Z8��Z�tɟQ�}���S��Q���a~U_�X���3s�ĚR]�$�fh��ч~k��̮G�jX(؍!��O��SA*_�	��Z��ExpA��Bu�+q��9����N���!��i�P���6��Z�t,V����\<�QO\��0�3�q���2A1Z��UY2�߁�JQ<�����l �d��.�Zo���tS�h3�vc����Q�v��l=�)���d�U<�tr�Tk��@�^�q������-q��=A�zݟ�b>�l?Ȁ� V��/��f\����Ϲ�.7w�[�#�X�l8��(�Z�����7���=�X� �2o�bQ�4�D~��Y4�{}���_�:E���Yb�掽�"l�?ź~��'�-%�u3}�F�]dD�[���`l#�ڥ����\�{C�����k��)�%Ǣ��RZ�S-���W���Hej�7(����D	R��-v(x�8�� O����R�v� K}���0γ�aU;�dat?����ɲ�yl���v��K]�-c� Ji�"���W[vS��COH��[���.[!"��O`z�q�3*�}�W����4	f?Lv��v��ofߗρ"�j,������l�T�ZC4�C�����sH8���u�m�l��)n�E�:lcWz��OyK���K��+l}��|�O4�0@a��B,�r����Gs^B��VC<��V6�Z�g�:�,�~�X��e��b%�+���>��-l�����|���,!�����?�i����>gνUP�����fl�r�K���/\+w�+'A���m��3�B�����!����-|�e"�7�]>���S���W_�"Uz�����<�p��#5iñɃ�=Lмn��v�{_I��	�r�S]`2�dSS?�k�舠?�.		��*:8�<j����j�������'���z��q`_��u��Fc���Y��?�B���wAO��d��UZ��60u���f%��x!D��#�{���R��Pb�hR|n�����q!d~�P��Mt�`�H�H�K*��<j�P�����`�����乱�V2�W��;D���9�!��;�m\V�g��V;׷\gW=��n"xi��!M����do�Ǐz��������#�b���7._z��̏<����I���U+����G�n�CV)�s6jwV9
�ढ़)ߌqF�Y���'2���bܴ�}G����mL�	ϩ�|�I���#Ny�+�T\�$��&�K����s�V��w�ؾYEF��-=��[�UW�+��hƍ�U���xa cJ���(K�mT�.��B����
�����r{�3���͆!c-��	�l�b��ڈ�X��N��.:%��GR�i����It`�A��uo?nF���^���e�;��_��A�xX|���L�7���sk�捿75��*�CL.;^�M1�QL�ʘ�� �5�Q�zcչ6��
/���E^߳�G,&���N�P =�Ot�`��Kbr�,�ɶc]C��9�kA6�NH'𬡱 ��؟�<�Ƞ���K�#G:�&
Y���$�=?�<�>��hH߿-L��j�$e���ݧ#2P�����ժ�z׬����c���L��6B�b?ͤ�bFx��:����&�aX�q%
�s��R�/��@����-���!��������h !��~85F
\���=x���_�v�C�D3D�I'���q=�_�F�ѵx��n�4't^��h�u�%F�q?��S
�xU���s�:�/^����Ͳm�b��K�š0�&4�a��D�G��%&�S}l6KbCx������uS��$a�	��ڿ���^���x��kr�\������|��Pa������U�mN'ޝ���A���C����6�5P<�kPm�.	�Kj�J��qXZk���#8
�G�h�}�7��X/��њ��z7s)�8�8z�W .�6��C͹�8u�-�G�<'K�ϒ@��)͚��N�����#wy��G�Yʪ����tW�d\y�����/x�d�%'yJ����Mp�v��2�	�A�;x�N	��߹.��ɨ\,zh������{��n_��a�+�[FT����o�J���D����[�[X7�x7�V3@.T��ԴI�#"���/���Bq��-EI�x�s/ys\�Z��?�hK�����X��.Nr���}�YN
2\_����9y8ZK���~�A,��M'�w��F�F[��,kB}� Z7*��G;�j�^���{����\}���yGx��� �Q2J"�/H`�d��=��|�� ػ!�w:Qń	�@z�Kٯ՛j�|�
�Oa�����a-�~�3`a0��2��^��B-B�<dk4_ꖕ�g	ejDn=�#*�8�D�@UT�׼/�^d3VplI�J:<�Q�Y8�;�*}B�5-�^M��­�iA2�UÏ��O�=�\�U�Kc�XK����D�]xE�����W�)	�c^M��p���N��d�$��#+��9ݠ��C+��\�*YR�)+��G_���1�L!��j�a�<ם�� OT�v:�6ȷ�-�z=�((�E2JU;�*��ߊ+� �p�7sOUaۼ�>D�;��k!��Y�����U�c�b�	�%x�u�W��6���z��id�l�&f�	��T8<�y0Zٴs#qK��$*q���G�C`:�8%�r��O`���]��1;Ѵ�L�Z"�0`f��c"��*~O]l����ƨ��=L�N�%&A������j�n��=$Z���*�,������\/V��D���ԐQ$6.v�sr#N�Ò���~:?N��04�ֺz�У�^YFN�伙�}��=��c�rL��x�م����k3m�/-�X�/R[7�Zّ���"%�?Oz�?M�P�e4�W��K�}������ʜ�9�k:�3(0N��@��
���vWl5�%�l���t�����kW��x<�求+�	�C�����$R�+��É��̠#����˸�~0;�q��FH��}ӳ��_�L��i�GT�C���B����r��Ϳ?��,P(��t����<	����߈��<KWYl*?io�:*U��	Ҏz�9lB׺��8;z�$y-��D�QC������?�J5�	Wk�bcz�vi� n Jm�D�J,���k��z����d����}�>��UY�������:�>F��&^��7-�8�lL��`�|0 O/�S�����<�s��ao�	h�z��uA��t�O[{�pF�(��ڻ���S��>S��+���\��#A����V�/ ��)s��̠R��N�O���&�VTqp�wY.}�(�D�j�/ƅ#9�<�[��>�ǽÎ��G��a����? 4������b�K�6�\��@���Xٓ����;�ܤ�p慹)����e���5��W�T��g�M��D��Z�N�[���K����\��H�7��`T��y.�8���Mi��=�E���D�88� �΁_��P�wA���R)oe������y���{����l�
�L���p�s�]�
��>|b�H�� ��]���:p���x���ꘗJI&���p�s'#U&/MgD%��E��w�;Q���p�h%�" ����uo�A-Ţ�G��"��T����1��lH+�h�����\��oZ"t���1[�����:�b���E�k�X�,��	U�y[��Y�P~��1N�֕��� zP5%c��=�NOO'�Pt� `�K܀�8�9�z���๦a�ixu�,9VW{�Q8�G��9�f�� @��b�����J��	�Ў'-Cn�,��c�V�V�L�;�@�A�1f)⵭�(_���I�`{ʹ��ڀF�ϕb=�ػ���b���Ƴ�s���cH�u��YY�mqL�������1Ez.�U�|������A@��Cٌ��)<���!��` ����5ӆq���U"���`��LE�����՘ʚ��5��̳��6\���q��l#Q6��S����X�æ�P�ևM��*�z�@cG��t���.=�G����d_�Z�x�x����ɅYn��}.�xg���$5��\�[��M4sܜ��Y��#��>Ƌu�N��	���ǆ�1y֣�u��>�\g�3���jX��qc��$[;t��7��m���ϰe���ˈ�B�zƥ�LS��m,H2��]J�:�7,�`��^�e����?�YQJ���X�%�0X��+V��h�-�Ҟk֮�EhnD�u���oĭl6/8�-t&���}��S|E�!������'&�h �ֲЯJ��O5�-�Iw:>~t��xi���s��:���7���=]����g��t�	�g�|n�<k�g��|fz>�v�����i�&-�b�KN ��i��x0������v�QkЄ(�(�Wo�v2�g�<����=E=���IU����ť�:1�U�������j�3�׷��`N��/���(iQ�9����n�z⎻��W��t���z�\���Ł���Uꀲ��7���:x��ʉ3�OgH�6��t������)
M�|�f5S�B$�����@LÂnuru" .rv��`�2,A��@��_�I�Z����� ���JxF�<N�A�q XH �����A����H��Ҟ���[iQ�� �!�Q�qf[ڪ4����!�Џ����5��o���rc���qt��q4��]m��is]�{\\�-�K��F�7W�T(yl�A,�ץ���u��8��d�}S�C�}�Jv��0��AK��sџ��@УW�5��'��=$#����}���w�$��L\S�������j��y�YfࡻxS^j�{�+Ֆ�6��E�9H�x�a�i��nq��l�C����N9��(��1x�oRȏ^x'�Xn�N���l�H��/�h�pO�]>!Ͳ����B�̤�|��Q)��v���!�ɜI���Y[�ᛡ�v��P"OW��Z���v���;�(����]뎂�?1i�o�+�
A@���u��V&l������үQ��c36�*�=��C��<��p�8�h�f�a�k��#�g�_3w��Ϭ���H�2㑖^RԿ�B8���8�ڧ��>8XX��p�̕$��Vj����	�m���/�^�V����Z�/������q푒�t�.\<�F��s�Z�KE�L1�ɍ����(Ә�&V���Z�'�^XÓ������.m0K�쯌X�Ez��\*DS�\j����l\�;v�D�f(�Q�UڴUk���By���n�6����NǀcfM��G9#�8��B���J�{P�D�o_����T�1Β�H�0'Ң��c�/����	�j%O�;��v$Nh�(��9��D�����5��5� ?�Ӝf?D��5'���M/'m�|���!�.�5��u����[�	�)|if���-��%�J=��l���9J�:<�گ=*�DuY�"�ˁW�H�?��+�c���$��(A�F�P���Tt2W�C�
F��,k8���U��˦�R�]�~�@t�5��B���.y���� [Sz%&��|ڲZ���|i#�Ԩ�ۅ\#�l��e6�y�~ǒ6���!�E�M�'lD���j����v2�I|Tz����0	�Ϻ)v�Yk���E4ݠ�gh"o�KK� ��<�FoN���AnBMK�W�����p$�<*DX>A��ͥꐧGek�҉�c�24^Rd"��8�?�_��'moOձ1�۰�g�t��~�u�
�q�L��\n�1�Zce0�PU��sZщ��0�>��1d��8��Iդ�%��'�KyjK��r�Ȟ"�ۚ��ER�ꨒ-l.b��b���s:~���
�dϐ���;���R�
{�N.�Ιj�����,(*��'2�:�m���i�ŗ�SC+'����L���4b9�=��)���{��@-ď��[�(�,.������Id�W�*�= �)���n�`�