��/  ���a��|[�{-r�#nl[m�v�{5��7MZ�|b��}�"�8LX��(�Z�ʱO�'�Z�i�%��7�B�^��8$�0������P�5#�E��w�9�@�\V1����,��r\��>!���N,��
po�I�;ط�&[��� �AuxN������!^�0d��o߹���ɯyw:=G�`�9�PyCE��8%X�7	]�*����pogU��(~X� ��Vrv����P�Uh:l���V�	�$���p�2��_1y�ȯ�u� 4�D�M��hݿDI� 6�pn�l�!`' ��-1�=<H_6�n������8��Z��,[��f��x�j����`�뻪{�~�!ټ�wF�ȉ'����jd"��H�X��]!�NAk!n}_��n�90u�7�;���HƝ��oN��t�Ҧ�E����U¬ӳ�a�j���}*8ʘ�
������@���)y�����	=��p���i*D^�g��i��@F�^�b<��?����W�b���jЦy�����1��������z`�J~��r[�Q&H(*��ٯ���:~�)(g(&����"Ƚ��.����
[�b�ox�r�f�:��s��a@^�I�#=��b���î�'p@�t�x=/��09���+�s�����-�J<���։(���ZI�j�t���Zb�f-&�>1b݋L�Q�7�	�;�byi���K���?F�願=̳��~k���I�!j=�m�{B�#��@.��j�e
#�|;�ꠅ;�HԂ:j���������=,g�ĵ2m�j���Pr��#mh�b;kɾ\/>�Ux�!ؙ��	�ZZ�-[�9ux�*�P�kB�M�� ��HW,L����nt��h��&���,~6빋d�i.���#�b���)��D�H/�7��z��ub�-� �t:�[�Z7�P���oɶ)g�M=2	��*���ק��%�����4����#mi��L�p�1��Z������.�e�m�z�z���ZA׈Y��g���O����P��!d��(΀�H�7{���Y}�\�����4��7,]܉
:�e:5^�I)y�`��R��k0���G=�-=�����[M��h�'�qC�°���Mp� ��ɜ)r���od�X���c{�������#1��D���Uj�����ҬxP��v�j���KwX-���3�9�!���A-�V]����	�P$�z�XZ.�w^y-����s�+��C�����D-�7��c�bE���ȅÈ�}>���7Ē�	������H��I�S�~��f�BA׶6 �Y�]����<�z�ä�����-�ʎ=W��<};�xU{�����G90П>����m�X��XA���OQk�;����-,� �*(d$�w��9M�[Xp�OV:�2���Lȃ 
/y4��yj���G�xソ�� Ê	��_�7GV@���Ksx{��n/1���VsÆ>�QS���&��ΰ�xT��]���'�b,��;�c��L��C$�|��nt�e�y$�_\�����:�!.T�[�E怦��z瓩�h�������ڢ-xd:36�^ѻ�!�/~/����W
���.E�h06�������K����+پ�|��:V�|(�� �� q>�m�G����9��|���m�e�X�� yl���ɺ��םX�RW���g������.���SiC���s�\�ފ֟�dB`���8���I֧��3]c��ʼ<���o|�+�n�n�-5�v�|�.���Ԥc�-8�4�.g�YNmcr�׶1����.n�{h>~g|�KN!%C�0�C��I�l_y���!�T_�%�JN7�FQ3c'̿",�!ܢ2�#�៲��`��(��Y��B��\�r�K���,�<���zEN�� j#7�ٶrˌz�p��y��ۣ|h��[�&;"��Y�&A95�K��n�F��ר�E�ĕ�<$oŷm���|&�2Y��6��rV�R�G.�<�u�3��dՕ�d�q�x������t<:s��/�ӷ�~����k��$�'s;�Ӊ��r&D�����Ǳ��� T�u��t[�'�Ɲ������}���b�������clh\�U���?zz�%��9�3�D����,X�g>_��'���ϥ���Ө�TM�}n4�d��8`�]�u�Mڷ�H�-��V��Fd�a��cdP
?��QKK掗H���)��JW�^�g�w���]�/P�����x�A�{��T�4L�.�3��k-%U,������!���1gvկ�ZK"�9u�k:w#%�u�d�X7�q����_T���J=O����|u�D^>Di�����ݰ������dנgņ��b�7������"�jP��X���\3��J����f�!��
���j���	r[Uދ�V�G1њl� : ";HHn�m�h-ٝ h��|�$�;�:�~�܀���P�W��a�6JI Nx�0Y�CMa���]x?"N4�fT��&Z�y#L��Kɨ�&l�����f+O<%#��t�