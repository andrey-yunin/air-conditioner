��/  �����Z��!=�.��$n����Jc��R���|4Fo�a���m��<\�\"�e�jj`�)�2��8T&����pM�5�L��-F�Y��D0���ݬD����\��$��z4AE7)�n)�,%���*�'s6s{��q�t��I�}���t�LC�:-��(���!^�0d��o߹���ɯyw:=G�`�9�PyCE��8%X�7	]�*����pogU��(~X� ��Vrv����P�Uh:l���V�	�$���p�2��_1y�ȯ�u� 4�D�M��hݿDI� 6�pn�l�!`' ��-1�=<H_6�n����3V|ߘ+�Ǟ˖���Օ�;5�������=�� �a$∫�1�S�fjZ6���`J�D�*ZU�����f+�X�a	P�1;�T\�IX�\�[/�y#-��~9W����J��~1,�����r��/���.
�Z�1��5��A����C"�|�=����ᾳgu]���g�)��׉f*6��e@V�=�x����`bk���I�ĶI�Ɂ� ����~*C��0l矛�Q����n��sM������ �q�0�4X�wG��CPA�{�@�g��Jz����S}�K�~��ˀ+�k�52c���\/kή��+}%��&�D���
��6v[ ܚ�'����%̗j�l����r��iR��ʎ�(�? �ac]7 ���Y n�&��z����¶-�4��e��Q2m%�6
�g+����M$�U!�Hl�7�p����>z�$�T���4��)�0��0��Fֻ��C<�y°��$C`�G����_^�� �'+��"�E�����~��B���J�S�-�ș�kP� �����]�:y0��&S55�ku�D����4o�(9K��,����ުa�*���8?	��+19{�&B��r��fCT\s��P�}&�D琨@���7H����ieKO0>�U�i�0��b$\̝�lRv���=���n����t�/�����۬�irӻ'����HL\ےeE�|����d�PIk4�;���.c�A���F���v{oֺ!�E��qW\�9�����sQE3MlQ4q[��������{��gjd}�.{�<��$?�Z���j��4�2+ma�Nu��,�f�_����E\R�tfP!�!���Ol��i"�G��]/I�~v^U xw��t͓�H��a�?7�s��9����`�]=4	:�Ƕv�:*y�,�p?v_��3X�T��Rh��\�d��ʱ�kǥ�S�Y���Ds�o��R���܍�]�ץ�JBY0�Ɉ����q�'�;�k�����'g�vGw$u�cM't�+^�����g#T����Y�$��u^X=3��*�����iS�&�eN�),H�������`�}r��C�����'���Dc���,@'�^/-2��m�̫uW�xt\����ͣsy��%��&0*S��WM��!�Pd�l2�M:k2o����%p-�U$����6�ݚ�<� Auy�8,`bֹ��r���} eW��0� �8����TZ>E�V5��~SßҐ���g�|)ǖ6o�d��.���&�=�t�|IC�o���c�ѱ�Y|����KiQ�� ��&'4 2��EKg$n��j�y�R2&,��Dj"�bH���Y�v?AgP�!j|AA�$I�s�A�"��I�17�|�79,A��B��Q]���e�V�;N��s}g&(=�w2[!Ϣ�+��U��c!^
ǵ�L��Ҷ ��cǗ�D��mA���� ��l�m̽�v�cE6�\�Dǯ9q�|WJ.Y� �j����G�hL�i�#�oO�:�T���~�s�s�2��N&��8�ue�q{�'��F�^��lτ�\9d�3�u��S[^ ��pǐ�����2>�Ư��E���%��0v)�}ʇ\by'<�'ЦX�I���R@�'>ñϚ- ���\~�s-��~��8��䌧ˆ��f��㇆{O�	�e_�*�������>�*�}$�F��dA?�q@�F�ۙ���:Z�?�+j�r���i�M��Kg�4��s��-���O�����I�xF�[�wOw�,�Z��"����#(Y$�op0��3s��Ɨ����oP�������(o�f���F����n�������nn��c����&߿T3|7U����dպ`�7������1��ħ���jo�v���j���\;�Μ`Y��xWxU��^�8�/�������*L�L�7#-aqW�E畿�_��.m�?��w	���]B�f�Jt�����V�.�e�^�AԦ�q�2-I�&��7��>����DSg�ޅ��\�k�8(�!n���̲H��C���뺀'o;i�Er� �C�R3�>����� h�sNh�VD��?��*�w浧o�d��&�:r�1�_���u���l�!�x�6�5Ce��̉�
>�^���c� ����i�2�{s��G�(8���z����Uͣ�U�H,'�#�ݷ�N ���gN �b@�d�D��������|����7h�@��,-xjF�z��8�nO�d{���V]Md^�ht��9ˆ:nR !p�GQ@�B}S�fH!V{`��!Uc`*ɽ�/<��bU_V�w��Ҽ�SU@��Z�@��馢�F]�7���U姅}� �&|?��5Y]��!GÁ{�(U]#�,Ï���1��~�G��·<�o$��] <i�q.���v~�
v�IΜ�����MT"���Ro�����hk����w#� �g6g;>�#^K�E4F���ǐ?���Ѹ\��0�r�W��{�f&<�gT� �������)]�t�s~�B3�+�	�a�W����)V��+qɬ���zt�T���fR~}��k���w�ר�s���.sΚ��H�^aȃ�.��c��5r�~ˊ4G[H�YxuQ@�R��,�&c2�=)�ܧM=��׭lXb(N2v���,	c�ݫ����fǩH,{�o��q��^Y��e��\,����:�=������~e�ˬ�p^YU.ehC kw�i�Bb�#!k����"��d~8�k��)/ٍ��~�y��N���Obz3��qF��G�^Ӵ��ce��*���I������3_�v\u�~�b�Y_����:�8�����YHZM5{Wn;��*\�^���뿗���C�+�$TP�/cH��N^!����CZ���n�s��Ɏ�4&�mn$��Z���䄛�RZ�Z�$_p�!]]%�Y$J'�=4�e����0�w��J�-e��<��B�� q�[#IFˈK<�Iu�!�,���?m5?�S��e �^5��C��I�}rB/TEͷ��h�$5�ZH��\�9�O�x댇�o_#�*�dr�Ԑ�f�	��>l�:F�r�����Z:Dzl�=D�bXOm��T0Z��+��\�z,�KL���궫Q�s�<�s$�y����w�I�`>d�k�Z���v�_���+�?5E��:r	"�OA;Ej\�s,��,zQ�~����uw��a1���N�DE6S���։ȳجBZ��[��6�����vW��C��jITƙ�5�f�KM��&�Xyv�G��EI�k��%��M͸���5*IF�W Yf2���`"��M\����%�� f����m��8�S~D�ޏ2�������aR	�>����px�9����������H��U�{��=�yĬ����]���2
kN����eH�O�x
<l�X�ɤ[���4��Z-������I���ŧtOw4��b3��5H���PEǱ��5�������,LO`�pY�R�G��������Ԙ�;�����xB<���A0��C�E���O����F��ٖ��~�d�1$���3#"�!�^\��(�r�(�z�O;��&E�>��Q-~���f�"M�x�� ���S`��Mv�r�g��Á������,W���:o~�� �e��{Ƭ��S�h�i�>���kt�:?#�l��%�"��2�%�&�����f��ZČ�)�R�Ч��d����^D��CG+@B%� ����j��_X�q�%>���بVXF�3.�n;чm�xǖ,��r@L�k���,�[����BM\No�����ăP�1�n8��H�7�4��{naCƭt�Q���{ȱ�B+	�B��q�e〲�r�� �˹?^�7f2���v����Scɘ�
Or˝4s�����!DG�����h�!��֣��ӳ�O�;�׺�l����g�E�Z*���U�=td[׿Gǻ�@{��W�񟻏;��`�x������j$B�-�<�?v�&�ap�0�#�)!e� ������S/L��qs���e�77�{?a$)&ܷ0pO��ܴV��_�����@�ܙ�i]���󗙏��dXM�F���O�!�R7��H4m�Iڪ�����~�*�$��x��D�_�
���g��� �}c���z$���`��L�ķ	;{}&~K���Y`S�*<`[�^,�zzc+n	T�ü	ܛ��u@��m~�W�Fه/�Mߑ6�/a%lSf�ٔ	�6.���X0���7r�z��.�N���RG���P�����=�,���
��Vq�rW�i�I��B�`��"�I���WZ����W@�J4��*y�^��]5�"�e����|�{�%8W��a*)۞P5�i�9`��S�n���9K�Pk����fJ�Z��u?�싆[�4��N�0i�����wuy�{���GA��ҩw��lF�	�G^�$���Ǚ��Ѷ�	��sJ�s�Po�;�ɳ+\��#��z(R�� =3o�H}��NZW^*����޺�E�U�Uy���߽?l���$�L�t=Xf��,�xDw�ȖΡ��|��%�v���/�:��H��I���!Ѫ�Ÿ�&�2����W<��̬&���%�&"d�5-�:�s�-��1]2�� ʿ�m��"�@HQ,��ޙ�Pnz��C����q�@vWҺ;*�
�M&��������-���'�˖$D��y��.;r��&�~�C��P�0X�1ڒ��\�T�)�o��t��e��:G�ԗ�ܢ�	�~CL���x��/�����yQ~��0�|Bj�������έ� ȅo�o��>�Ll�5fol�h�\(��*�)Y�I�����š�G�.�;�W��ߋFK�fu9n5�Y�{�@�W*���s!�3'9c�����M{�pёM�ISP��v��������Gi��dq)�.b&=�lR���g���VoM:��S.V����vZzr<�l��(�ʫ�q�iv'�����^Ϭ��ixxh�S���ՅA��	��1ݰO7�֛�?<O0/5�؅R�Wfu�������讔j�B�lq�c���:�'X:���h�0,4�y�Ǹ�j�m��_��\0bN��K9��x�ne���U���U�Po���Q��_��p�}� �8�1%�ͅLz@�l� �5{P�Jv	!��yfٌ�'�|6 ��$�C�N��9کi��X��̉�����w#w$� �%F�})��'Ɗp���8^���K�'�i��chO�>H�9�[��O>$�����6m�����9��t����`�m�����VϮ�STǿ���#��4� b�YF�N����o��4��|U=���\M����k�Uʠ������y�k|���A���8�� 뢄+j�}0Y��"D);��ԭ��i���c2y��%�@�T�
%8�°WZ�>�	�rF�S���:��J]F�F��#�T���<��:C��@N���2����"�j�/ǘ������)�n�����ey;߮iC��\߳=���E�d�<�5��'�o`_��`��`�Xp!y�B�d�������.6@�=�j�g�)i0z�}�� �����s*,h<����<Cmɲ �Iѵ����i� ,Ӵs��݌�~��Ɉ{����6���ڝá��偸���#y���遧�W�lB��\ӡ���b����t�n&���<�n�|%�C/n��A[�;"���n�Gbh�$��&�m^9l�XbE�l&���K~ ��c�%�����%�f��T�9�m�V˵��"�*b�p��!�m�;�6��'�ί���YTmM��P}�Tx�5#:�LG5P���V�Ovq�*�kp��ßA�A(���tV=t������N=ݙv�JӜm_+�=>a2�2ȊV�O�J�
C�#���Z��W�j�G�ghɌ��s�  ��٠�ͦ���Ͳ1��U�jBh��Q�S�5���tS�sF3� F���
�Ta~��	×W����Fb 8b�ב�[b=1o&��F���J�������3�D��D�Ȗ�Jbd!h�4�#}�ѩZd�����&,��#��r�BX�;�G��8���ST���g�Q��ɐD���[mŇ�;����:�g�
t^ی�U05�6��� ��9���.�X�����_�������2���)�4�D�$�at;��Q&�0��j�~����hZg�j�������T��\�9�j��L��"C�]�pi�����&j�B�&C����3HA�M��l^"������������*�B��H{�=Γ=с7��D��)�'�1�qEd���*QC�d�1����{�y����o����s�����*��/x��p+_-�V;{/ݘ��^���,R�1�&U����H�IiY.��7�WM�+�U���>AϛE�V^I�iM$�{Fym�6�#�1&��HD�7���q������T3�2-{X�]{Kc)�]�|,)����*A�T�����W�÷�Nj���:�@nÑn�g��C��ҳ��MX�&o�;Er�@�f��!�����ʵx��V�0_�͵?���̤%)�UZ�o�{����ܙ�X��L�O)�i9n��c��a��Ƣ6*+�=�jq(�iu�K��d,��Dw)E�'�)�H[��jSO��H���>ne�����jY���[5j����,�� }��,PG>Kx��g�c���A��+�\ŋ;uf��	��z�R�#^�Ɓ��>0o�T�/�[�  ��&2�	s�xT�������8}��$�y��Glx)9��^�b��<,sXk��?{��^cre�8$�b�>cP��D��.� �_��uQ�ER����}��M�-�ָ�����Yi��nv������<e�Z���}�G[ �.�s�K�|�'ʕ%xh��DmX7㉒�sz�[��R ��(�H�u!�z�B�$+ 0��$R�e�(����#��SSl��Q�#���y:_����1![��V�K��t�����t΅�D��ؙ�zd�-t^�ۚ6E�Xk�M���R�DC8.�ۿ�r� ������ѲZ����sH�"`I״��&���r�%�<��Lɴ@���{u�<����<��Y Vȡ���b��Ϡc�Kд��>�m�٦C?�73�yc���޹�9����d�MY T�o2{~Im,1�1�Ƀђ�4l�~h��P~��w��t/�K�v.����~��2���$���"�����KsD�����ݓ�؍
? �ex���r9���9f.3���4����OܞwƄ�}�>.͚cʠ��r��-+)>��7��HO�o�aK�.�粅&(�#)�g��6�oj�Yj4?k����?��aS�Pܴ_���a9�9bhry�@OLl�qO�0���nԿ�z��9s�,oß$��5���#O�z����{���J��k�t�TW;�N߅Y	�߭��{�[ӞK� �0�H����tG�o�c˺o̜Z�t�U�P������3��(���60�ozh��z�E��?6l̴!�N#ڢuu��wş�խA1�������)F�xXCV+�4�kx����0"{�3��tj�&���)�^�IyЯ�� ���@1�T{�QɅEB��|��+����CT�`K���������e��@��J��{H�h�L�X8�s�񸌬���cBo��!�� ҃�&}�<��lӬ�i�T��!"Ƈ[�9��L|���+w�v���� �^��5��yE�w^`8&=?)����ap�(u�G޽A��O��>��`�+�ZR����c4Mw������K�+8��K��<����rFsa-�n��>]|���RE��`PAsYv5����9�O>ܲ6�S��
�9L�=�d5���u�!�{+Ψ��iL�Uhy�u���1f{�y�=��=��!�7Ci�[�O�o~��y/<I?�v��$S3���jo�G���z~&��谚�9��($��۬�X��Y�07<3]~$����@t�{�Ǆj�|Y:� �$	c�p�����r��
Sz��s��� 4]����t�jd�G���L����ir�ҏZC��9]����pFlt�^��t\�Q*���5��ż��`.1�Ċ��3hFG�buP���d�T0&���(��yt���bᢜfqDǾU_�V�>ӥ!�T;O,��¿D�؋̑���2c��ROVm��G]௎�v��&�'Xt�alpC|�H���>Y��oF@�g��>P���&a�qAsu��R+<�yy��2�`�]�<{Zjq̆<s�p�dR+~P��m�.����OGe.�īd9|��-1�8N�6�a���C9��������O��J�1,�F��O�~��-G�O����<|&6�����K�6���6x���~n+�;�a���XLX�k�|E;C�R��f{W}X�"8>z|sI�:z�V�q��" �]_����O(��G�a�����"}��ui���.3�ht�6�<���G�������MԽ��R����B�4�w^>8�jĘu����_�A���"�Ȭ���t�B�ed�/cpƤ~��4[�Qnd[h�	^s�ل��+�Z�Ζ?�
�H��b��`���������I�_6�o�WO�H��*)��z�]�F�D�r��#~�j��`9'��Xz�X�)�F�t���,;���K���}/ä��:��?/�q����f'���:�aMK���k�$�0ey��<�� ��>MGЧ���9x5fm���Ďk��Y@��`����W�u�R��Gzuk#Y6��d��WZ/W�Y�0��"���9C�(��O�ò�kxu3�EPL>�3f���F�j^#��Ur�k|M��tG�XĐ��p�ua����"M����
��ё�iRB(��T��u��M(�e��ǀN*�ʳ�#R^Jxg�气���褆7�����+J��v����p_����;������D�]�ϴc���'
�-_G_Y��=�<;ODB�������	�c$�6���7M����B�[��=��h�W��,T�>_4IN��^��������X(4�����#$��T^�'�@�W��ڟ
RL�`����@��k��[�0'V�� ��b�^7`� 4�n�wl���,8g- ~�s�3�=G:�0���bN �2���m�.OWK��z�;'�"hE+�kj),�z~� J$Dt/?��(�(�VGUW��;9"ƪf��^$º&��*ky���(<b��d�#��D7׎I�P�H�n�6I�c3��l�|�Ή&	��^���g�Ow���\�rh�ԯ$XD�����Ǫ�5T$�k:2/x�`�L���A��P¹_��W
?oܵ�0eti��EוB���+a]�+�̧�	>��x��G��7��������T:�;��b;�zS��>��'���~��M��q�-+,�A�J7"��VH\��0�VJg@���0zR�	���4���A�bֹ���_Nפ�=s%B@�.S��Nwn���CC�,�x�t
�#b���Ee�����z��b�B;�B�x�#ס#:&K."Z7�])Ɩ�a���aPGWå�K`U���������Yq�����$ ��%xD@��D�#HP�q�R�0��(`r��q�a.h��!"��U��G������nd�$���J��%/d̢_�
A�SD���v��\7�j2��<����쿳���v�b3�X��?��2&C趐)�	ե��]��#��-��}���f�Y7�_�prX����E�F���/�-o/�"��$[� ����*����T�)�����M~M6�ܘ�r����d1�5����V�l4�E�ٚ��b���S�l7AkMn��qkF���.�n%�������b,LnHT�4��L���7�!ݑ��T��]6`����P��#�g�k�U�Ɋ��-�DN��aj%�Ӎ{~X2�B�{�մt��e�E������U���$;U�13���R�W��
ߐH:R�:h����'%��)�vN���Q� 'M��KB�es�LQ��O��<�rS�GǊ=�~�;�Fș�6x�2e���MW9&Po�F��a�3^�{��X*�ra����m�8��ۊp�*��^�Ws�s�ǀ�� /�K#5��ȥ*�v�6�	�����AL�#����*�����w�!����B�*p2�)X�����8î��X�������FWN�'�6+OO����`�D5W��*YU�#q�k�7D��b2M����C�0�7,��Ӎ%�e� W���̻o�LN+U�m���%�.�	���.��Jd+�&��9X�}蒆��f��V�����}��珔a���.3��o�Y��8�ZT��c�縡p�uǄ�7�,�M��Zz�G#�ՐZ!*����k/N��O7��o��O|��y� ����x�fy����0�TG��/H2N|��T\h~g�:��ƛ{j-�X�?NX���&�NX�4�)<�@�^#�ڤ�H�'1#�28�C�:v~s�cpdŜ�	���[�z?c�y���!�{��e��'f�������ȴz~�$5����@v�B��2���H��� �@e�T����c��N�ב���_v]�o�Wyf�]DͤP�8�3��v� 4�-Y2��^���eB��#�)�PYdD�J�6�&��e���l
w���r&��A{�O���DK�Gh �؍���nM��b�gp2�f"Yq
���@+8��o[m�������o%�q�+�J,��J�4�y^F����v�s�_�$2��ً��X99�2"�NI6ڹ���d�Ǽ��-�E�H:O�ܻp�O�#6>�b0���>��e���㷢j��5t<g�����f����G�!����M�0�%�jQfW������6����	ݎg|�&�>��;�	 m�7��.��j�N�^R�wq�pk�^+� �/�CX /���\	��X�q��ф�_0kgf�4��X�4r��j�:TN�K���U�Xe5�^޸}A�%��;�(��X�MS"�Bw�t���*�Ƥ�dm�J�M�C�����4���hn����2a���9̠fV��2���ح0^i�v{�q~e��N?ת�[=(Z��0�8�Ǎ�I��b$�c��`���L�=�r���>Z�x�xwu�����1�b��!�.ap��a���8��Uny7�Yn,����{��,����3DWfL��Z���規ን���g�nq��+�����\�%�ns�2�@@U���w���L��s+gS�h�{�ԎCBƊ��qG��e��h��h�邗��m�F��wR��V5��^�
��a w}<4M[�R�ذ�Ke��� 	D���H�G���}��
`:�V��.����lD�e�w���6������ڿ��5��_���N�-�������b���~A�E�-�f:�F���$��%��5�
�^�,g�-�+j�eC�Z�ÿ8�>fTi_1�[�4��w����W��{^[��@\�Y�R�>�73���ٰ��j"y�z�ean�����Ž��Eͺ &��: ��	��>��D;��3�g�F����#bk�rb⏮�֯���Y��� 6$�2a7��`]���R��+	�m�>Š��B4�����(C_�.�\e �9P�[��Mr2K.�;�'��5D�&$g�RH��(��ks�� K);q�H2���K�^�����%-ƞB� �~��#؉�s^E�Ҥ"G�ڤ�JP�nD��i��evD�@��&I�W���A\M���ԭ}n^��n\��YE �f������So�$�I�&B����NYSı�s����4��i�Yq_Ǿ�C㫁���z�h�)���G	c=|�� �����\_>[�τ���a�W��w����8��i�_���ۜu��m��:����'A��[A �jA豨���?�:dgӞm#:�3��/������u�K�mx�]��9gm/�q���Ϟh��L�����z�*M�L�,��-����|��tߺ�y2�n|i�T镨sڭg����r�'x�Gs��^��6��qؙ�R��Ո�꯬����{2�\ǒ62�D�~��(:��+HI�!�"�2�Ak���UhK� ��@*y>��Qs���~�wy����T�p�����+��e�:K�4�e��`�d(�C�ݾ�o�r*N(�ϪHG�����7�]�������z�N�s2Ӡ���_��}�H��g����1�����)�.�����y b�d!F�m�;�*�[ ��?L��x��C�����<��>�c��;ty�~�����d�)��U�eH�(��Ӻ|�ON�܍�QE5|w��-{���:��˺��}z$��O���#��h~̴L~E�@����mRV���lq���FWm�90��VH���4G7�R�%����`�<��w~c��/΍�R�J�ٌ�!�G���+|o=�z2?�@�9��Q��&Kxe�Ӓ�u��F�ȴJ�� ��eq�pē�~�i/\�}���{ߜ��H|^)�L'.�S_���Ey� z&r�x����ew�w�_�u���܂�O��2)f���VAͽO�B,�(��~���zx\���7�|�o����������"оv!/�@�I����Tc�b��P���;��#J&z�M�M�,�|CÿiVt+W��9�H <��{7}���Z��&�
�L_��_����JW.;����`p�s/f�?��q>L��/�4����������?���G;W��2�"Yֱ������t��0���'�S;z\��>�9�m>jC�¦aR(�b�dոd���U|�nd����6�1�b�����z;��15��tۭǎ>	�U\.��pppqՌY����k�����e0a�V	��PA�<� դ�$/�Ag?=N�.�^�J޴�r��k��a�&玩ԓP�n|����<�h/��.����K?NB��������1lE@װ4��u�=�5�`]I�%�GhN^[���!�^g��l��B�_S��YԴ��ᶃח������^q��C7;)/��\�Cee��A=%J|8a��װlO�m��;BV�r)~��`�t��7�e}�8oLkN�RoL���|N��4z_��3��JH4Vi�p	鰞���Ύ�Ec,.�4`�� '�7����;�(6�&�l�)��xp=Jg���e�|����,X4���	������(�(pёF�Mf	��Ts��,��7�Z����x5�6X/Xk]P�,���z�#2]��������%�X�4��#GF����� %,#���� GɈQ���t����j}�rќ��������}�b������m�h�A��;2jv�&������Q��s8q=[��rL0�XV;�)����s(�n(X>s�ƫH�p�}��'��Y;}�a9��tm�\�}�O�&�cC���=��c3�$	R SnX5��{g\T���9�R?��c��]�S��}�S��m��P��z�D�ƶT���q�L��Z)�;�%�Ԯ�e	:�p�2�Z��u�MM���Ɛ�Al����p�	��툖���ј� nN!@]<ꤡj���0P"�"I( �-h��&����2k��Y��3vK�P��a�d.JC�Y�X�����d.^�&S��T�n�������[�%�qwTka��&G��[�}��ID�5T�8%�^������߶��2��fߍ%��2�1x.o=��]O%/ZN��`��6��5��vl�)N�v������a�^.����vσ2a�/+�T�Veg���=��:5["�a���#�Y�ъ��G�q8�� ���pyC��!�_>��V����GD"��p.�}��e��N�*��ȱ�9V��W˫s(�Z��󱪂�ܮo�b��O�G���I�m�����m���~ޮܹ�q��0W|z��T��R� ����r�I���5"]��0Df"�����^^Z�.��eH2�^}�a(���|q����
5.��avL䧤(�1��ǘ�܊i�gTw �O.zt�4�K���ǀ)��"�"�T�l!����mx$>���Z��K�1�����E��g*����Et�k�R��/������B���Z���s�;37g1�L�9�e���#�b��
�s's�_��Ψ�S!�'��ő~�8_�����e��2�@-��A�8f���H�$��V��".%��
r�6� �|ç� ���gA�f�v��;��q�k�2�$E��H!�� ��R~N���"��@�xWR.�"2������6���~|}����v�����6!�F�%�+Ԏ���������˫�oe����ȴ��g�g���*
�&ERMd���؝��X�:OD����8��V��@�?v D2�[f+S�2��	�����I��429S��>�q*̵x�E��OȀ�t�uݯ������Y�0!K񲤽"����t��� ��9�lO�`����n8�a�N�3'�-���b��\7�?���ÓT����qzM6�Di;��������	����c�2�x��
P��yP��Ak�jp墫gL��񈲞d��U߯(V�ޑ��/Z������*	��ۥ������I�`WB�lv�/��%��es�N쮬/V1��|B�q��h�cP\�Z� �6�7lf�i�GQ4[����	y��]�m}��q�E�o�K�N�c�lY��bf(K�W���Ԉ�?�X�����8b��>����@/@l��^ڮj��o�T��G��.�2���֮���H+kh\(����h��,p�l�/�1�Ӂ�'&������J���]�Πif���u#
>>;��u�jLV�_�����4;�9dS�@�w�2�Kb�'aVbF�'pӶZ�tiz�������FEA�#�ܞ�Z�,���߱d�@�ԂH7� E�����2�/rpmo�]4(�<2|�}��'i��,�����9?���O�$��Yn-�%�Aq4�lЅPMX�1
�l�"{�Qm`[�⃴�w���9dOD(��rAw��[��ЛZ
ы^���RYD7$����@CժS_���X���U��1|A��#�J��̨����Bܝ���,���Gn�$^ZZ�bPl�k��K�4�'꤬��+�q�������~��&�<��������[ɫ�1�3�_�3V���(�etfj�>����4eaŊ* nM�� U��I�Q�����d%"xz�`��-�`�ݼ�L�rN�P+%��|�oZ�=r>p�b�ɴ�ڲz���Dʌ�K��P��oh�=^;�p� ~�x��t�1���E�̥1��؇:.��>V��A�taw��8u�92Ҙ��>�QM�¬rX�0���0��6�j,��ߎނ��&�$�x-���z�G  ��[p1��:Ǒѕ��U�)1u��y�b�U&�'�_lV�E�f�9�;?�<�1�)����b��";4���zGϱ��<	����<jW`�R,Zt?V��r��Z�Hs���&̼�H��ϑ	�e��F \г�Ӭ����0�_O��*��]�na?����DIC��H�S�~F"l�3��џ���&6���vi�y?bV��B�У�ؼ��!x��3>�~�����&���$Su֓H���삜���q��k$t_��қ��D��~[SϠ+���)��q�=�v|���e�g�'��N��;X�y�-\�:|�K	��G�f-�hK��m�R)n�Kk���c����Xp�u���C�.�a�r� �ﲰ��ڴ|�,Jb$Zꚗ����k������
R���^����/�ܞ�S:Ԍ#dl(�4c��Gϓ�k b���ٖ��R����x��Mᙼ��Y�n�7�g�ru�e�p|�k��C~;����WB)�]#��Zb@�~���^k���$����[ J�v$���U�P(V�Y]��E���Wi�:�<3Q��ն�$R�F��;�]»�`���i�'z �H/j���,�o�Qѕ���<2�]%��F}�]*�#,��uTI��(c�x��������9�TE�;���k��9HF��濴#�Eǉv
���@ԩ����k��)w ���{-�e{�m����P�q{[��zwpM�j������'IC�2q�UQ�)fU�uz)I,6�>�p�6{�~�E���hɮgٽh���O9}�q��H���Ry�8V���UJk�f|ˈ%.�̸H5Qd�AO��5���&Hf^�S�1J�)>|!.O��G��*ċ�S�T�c���(�ȭ�6:�	���猄��d�[�ŕ�ⶑ�%2��Dc�hS��i�_�j\���3��U�P\��K-kp),W���S7�C��w�q8���(�Q�m�dѣ����B8{���p�Yai���w����v�颌3(H(n��ǩ�Pi�h2�����=��<�4D	�6�<��̠�!�3s`�<Xߙh}���vMUtčx*����a�����/`0]?������$��?)�8q��,��ڿ������J��r�ə�9�I��44q����6��!�4=Ӈ�Ǚ��3s�и��+��i��8<�� p���Ã�Sa�Ka�n������=�ϩo��>r:����&��Q��<���j�� ��Q���!ָ��1J_bh�B�T�R ������L#�H��u�����g�'����
MY�$Kp�h��#�����Iswpָ�����8+&U�7�)��� ~ߛ܎ޟ�u��P�KK`؄̘�zX�IV,�?:���P�>���Bzf�5Et1����y����9^�1��A�Sʾe���#��]
h�v�}�|����#���t,�vK�h�VQ��'#�WR���VI�qI�z�6�j�<�dZ##;�s%���B�V�:¦ikV��@Yv�(�f�2�J�)~]�2�B�޹?�V����R�� ��v�)�MV�^\�8����$��=�����p0�O/�����ݘQ���].j�~0���ҐxWL�Y�yڪ��I��F؛��X(r�0���E{aaS���R�_V8��t%��ks/ݠ���"=�b�t�����9z��`_Vr�w8�釳ޑ�ԡ���A�8������Z�X��I�!�Կ%ڞ�Cq�)ĪC:�8E�,�h�ލ8��?�k��K7K{p��!��֔�4c��`i������t��K��RX��^K`��<4.�HU����~D���2/�9L�s5������D%4�r	�o�vho��Gk�*�V$}��ת2<+푒6���-�2��MP������
����,+8��h�N��a�̡��y���<��kJ��,�m��d���hN*bz1�E+)�A�}��Ь��eR\w���*)�y�&�M���(Rͦ�>��xqiJ��Ǽ^�#���w��/���$6u�6��)a-��@�BY-��3t�#G�k�=�FlqHgo��Gs u�BѠi]�c��=��&ݓ���vc�Px#�8Wmc�	�'?�zf�CLTg���w�N��"��ͻ4����Uhv$vkD6��*#]ג~��?�+�T����s�U1Jd�)��q�Ӓ����np�TN���K�.�#�n����y9���P��^�����3*�%9�����aS���)� ��넓G�!~��!�3n4w��鋇�*3Nh?�x��&V�ޑG�����߅��չ)�E��aԜuss���}�	P��.���dO�#_��|�K����F-�y�뢂u!�-B-�cA}�ᗉ�R��c�������y逓�K���Iu��j������t���y��e�l��e�o'h�@���6��K�Έ��fj���2�nb�۩��NH�����Q�0N1�'H/�P� X���{�ά��4.�~��P�#��Sy�������heB8��`�����7y�i?X�1W���Aٸ����<��s�W	��;��kmx@�cG�.�%�_��O�r�^/Nk�*u�⓬xx��e���
>�����|���#��r�f���<vm.��eVD�ĈV��<0�6.��|�yc���gH�31�+ZN?�0	�׮����T�� ,�+%-��OG��R�{-�&�%rv��ʨ�|�Tgゅ�J��Bم`��H��xko�#�eW�-�0��*�}��<��Z|g.˓��Ix��0�Ϸ_󏨁�	�N����j0���]+�^�>�O�7ڵ�*�S�њ���T8����;�H�O8��9]z!n`�<�cE^�����'>����TU�s�z��;y�� >('�|}��X�b�I�&0)gII�k�%qf{��"�q�Mܟc鳘&�#��C��� �)�i����VoD���V 6�Q�$��ϝ_�v�a|Oل�ćђ.k��}KÐ�W\�!��[ud���Au�QSC~NH&w����+��3�P~��k�d�͍�%��>Epw��&���.���M%\j��P���YK�=SX�������b<��N��N)D��2��R���'��N���6�q/|��T	�{�[M��LoC���+�-6���f�kZӾ�A����<��5�nտCN9�\����%��L���G�>����3�h��!��.1m�gdV]Њ��V��7P�լ<*g�D4���
jٍx�?�m�F�r����O/x�������8*֨/,R��1s�_&g?b+Z��,������f+�f|>+���;@ÿ<�4����/��S/�QB����?�G���Y��e�v�}A�����Ũ�� �wN��op�O*�1 R��8?.MO9_p����4�]f{�`�g��6��\{PGdП���$e�Q
9�jsؗ�$���]kHJ@B`n���[��!?�I�&>�G��٥��g�]��[���m���]}��(��,�z_� �]�!�-�Z��D��:�Mΰ5ckIyy֟����#?��+�:$�=�Ø
!��\�+H��IQ���ÝZaG���h�G��6x��ѭ�����D�+��؁ڱox�c�G@�4�@-��S�ۤ�Mg�x��|d~��
�#U�83�i�j��[h�����{
��V��O����:���DR��O�)owz7���i��Ƿ=��$% �u��O�n��4�jȔ8Z(uiko8�}��Ϩ[ٸ����s��Q�^ �Q��4{vH��9�v����c߄�ϯ�׳�	pvG��gI��qY�;�<����Pab�B�5����Ź����k���m/X��U��)̍��X�ʝ~��7�qޫr ��b�TZz����Jv_!��AS9}��`*|WM�h��8j����.�+������}0V�;�J�����߄�I��/�-i�9	`�E��z��h!12�����F�H<�?���7'�������vTI��������p�xdKSv˞��i�׷��~/L�U��_AI�^�Bj�=l�v[^�W\}�CJ+a1q������3&s�p)9�s��L��K�*��/Shq�_��\!,��{B���4M�X���/&F�7�L0ѹ��==Lf�.8�)��}K/�8�ۿ1��A Z�6����S⛐�pc�~����?�95	8B���fCq��9�֮AF�U� @[Y���?�B��|�}{p�ͯ��)C�n�5M�o���N<n��?��f�uO9vˋ�����*i�	�ע�d%|��	�0$U2[h����^|�b�
��wjqf�� ���W��M�
�X��_�,���[�-���a�S�0���6kXz_{XXL4_���gO�3�������a��O��Y�:����}��6��p��]�8���Q+rLf�B�g�)I��?��w�핡@�I��л���u��r������Ɔ��� �_B�0�Ta�ً��ezܘ�S�3KӇ�W�2��B�H�!��=N�m�=���3=�`�~XA�Kͬ�\A���/�J ΘH`Ϸ��������Pm��l��G����lEv�N\��;Opb��BgFT�
*<�|�O	�:�r�l��8Q	�%Sj{&��}��窣펚F %�`5������E��l��i!B��;�7
������Q�a�����}����^p;f�A�������+��d��OA
�	��P
��K�81sֲ��Ǿ����5	��ܪՏH���ŕ.BJS��pj�s[����c+�Xb�y�:�����-s����գD�L��6�K��_����d�>�N$��W��w��v�S���uR���5���>Y鐹b�'E�!ØM�,��;6�&.�to1嬏/����{�eb(U����Q�bj�l��üx�C�"�

|&�)�l���Ҽ���`����l׭�Y7id��!n��BĿ!z����Z'K$s�-#���� �T]5$�r3^	q/��@:e�4�.wV#* �Gz��΋���c��iPe��������蝰��3�!Dh��h�Pg�1d�j���ɷ9D� `w�^Ȝ�5�����xq�������!��:ҚP7��ҿL$}�d�E�}���d��EГe7���-�0�<���m �L�q���:����#(2�u-��q�)�y�3Rmd<M';�(S�.�>#ي�B~_�O�XN�3^6���e�|�yvτ6�Vi����_ȑ8�V$%:��f��9}P�Wh0��@���B��l��L��wL��\P֔s� (�˸fd�w�_���7�&�4�6v9�@��^%Y��`.T��c&�$f�;2Q2��>f�>�G��c������(O-���M�����j�@g`���LUp
�	�#�h8�&Y���a�^hĿ`���B/�~S|Q�G_��*��4}|Ɉ�|�y�R�R�ru��_Eau2���!��UU��!#�ਨ��n�Ax[+xsW��� ��f'R?Af	�'�a-V��$&��W�n�2"C���XY����$	#��9�#+��#��>�0p�!u�\)��O��[�c�Tڨ��Y��pa~��#|JW�q/7.��v�0�l��w�<�g5�H��˾����u���*���3y̫a>�Z9bi7�r�>"�9��جf=�A����V>�eȃ��Ӳ!���͘<����蜭|7i�.*�wgg�,,iN|K�e%l� �΅��׈"u��}���5<�!#�.���5� ��%�?[Џ���jJ�Q�3N5��Y��O��݅
�zY�<@4��n*���/hc/�8	��%w�� ��U.o�����j1��Dϛ�J�L�c�J-6�����W�����<���>�0,!d���v�,QB�c�H^�zaW���j� ��&<#_SjVu[���P!�D3�-��xiN�X{	y+��/�t<�&w��/pF��n4��|H��)���,���i��xX8F����2�Q��m����9�AG���*��*#�ޞ�ql��K{��f�Į��m@d0�)=��� ����8��|)�iZ0)N�mw6C��m���[Q�V�;C�c��0o�ϣ�[����	9��i)��5eVq6�Mk��0G����y��B@���*�"]������� n2)�3����r�Q�]�=���n�Vm� ^���Hi�ɢA��uy?�ښ�}�Ծ��:��*�|�
�Y(����¿E��C����.|��<zRu&��Oc�Rq\sk�S̽�e'�p�3_q�O��$�
s�NA˩�����&�ݷmbLB��(
 �D9���w��ҝ�����G<�h�3|�f�L�3�7���>M��!y1��B}mԚƻR0œpQ���?-�����'0�פ���c���Ÿ@��=;�s�c�����B��3�^3	��a\YU�9XD$8����M��
Mz^�r{x�<�|$�2!9m}Ҩ( S �L$��1j8�L��rXحfBX���.��Uł�aZ6�q^� �S~f`Ӑ���] -9�(�3����)��}5sTr��x�8���G�/��+���ݻ�Rlc��͞��oYz{�j��m�ҿ��H&j��k�\!�G�F=���kkO��	�C���F��*%{H	�;��`.�ʳ�x�c���\c��]��n�C���A')��iVA���G2�È��Эt���b��PU<���DR��q}FDJ��Z�x��v�3�.H�1�W-�5��� ȧ��OfFR�)�j���C�R���P;NI-q�kmae�m�vs��V*���
.$�:�
U�k�w�"�za�j,5:����M�n�"���+1��~��H�./!t �́��m��&jj�WP�˙|�Q����'�+�͒��2��]۸/!��q���_��(; �j��7��F	�9�3�qC�B:8SF�>��S9���1nl0����CK�]	߳���պ������O'���e�W&,Y��<���R��U6E��Bc�h�>ʡ��E�M��լR����M!�}_�e֡jy=w@J�I�Jkڒ�n�<Ң��ֹ��
i\�gǔDl�����婕ͨ#ęlM�L�m��	�T���L������Z4W���)7y&�e�$�N�}m���&}���x~�x�$�Qi��m�R�^聮mG��r��r�g����p�x�r�mu3Y�a;B�Y� �ͣs����Q��IM���HAx�9��@{���:c|�;g{+J�'����c/���v9S��X�̏�fvg�Ӓ��d�9�/V?+�N5�m�f3J���@��u�ky��Y\�Μ�N2��G�W�4�*�S'��f�!�������[a\_�\���0�{���f��Y�oL~��[.Ub����71�1�[����7�۽ZE�0�)�	�
Rf�R�λUѵ"26T����H��)�t���1y"�4�d1���}{�k>�Ju�ņ�������ztɱ#M�[�Ϊ8$ῄ�$��y��LDr(Q:VJ�B�U+Qdco�a��� ��O:��d*���0�bc�Gd�P�������q�M�1)�j�p� �ͦ]V�:��^������Q֬����	XE��mv���t��t���3r�[���h��2�e����&o	Y��:����ŕ�f>�W���q%/���N�FI>��Y��ko����q'���US!��L:n伾��?�iMC���^ ( c���}m���Z@�v�EN%��j]+���>D2�J�$�VjUu�Q�,�7.C�\�@?�H�ʛ+z�UA�D�5Ֆ�'A����D`��*�����s2Yѿ��G�i��X��M�"?G�a�_�~;�����^�Ƕh�]F��+�@�SrZ)S$Ed�}�6���V6���>��)��6_b����4P0��쯔��������4⯙:��Jy_.W���o�ؘ�)dM[*��ӎHQR�O����l�q�a�qYj�U]F9%�H�&���G�]�$��Sq����GS����ɚx`;�"_`q��eH���+���.y�Q�h�9�9�e���J�r���cᬑ���p%�1)�qY	�����٩c;\F���yxB�o�I�Z�s��1�P^CG�a�e�S'�ն0�Ԋ��U?�f�yh��$�S�ā�̉��o����ŕ� ���.�J7�e�%@L��٥��[��`_F9Çd���|^�tq�6X��,�f���E�o<Z��K=C��U��z ��;�Dp�ƺ)p[4���*��,��$�!UZamUa�kg��NF�Lv�?n���~��|d�ǽȼ,��x>z���5E�<�K��ڡ����a���k���
3}X�2�m�
��L2�;��%{�[��}�Uɇ���\b]Bݮ-X�F盄�"� Qe'rḪ�ƻ7/6ppJ�Emp3�#h��Ԧ׻JC��d���Y�s�D��2���x]3�ه��4g�C�%�}.!�C�ԫ���b�T����`��
��-�y_�y!
囉`F�[�t�Rd���}����3ZW �i|7߲#B�Ԇ}��� ��ʛ�X�P�cGVe��?�P��^�5h�Lrx��>WT����z��Y�R2��F��������b�,�#��όHFת�e򭌱9���_ڤ���M]C��<���C�yo�[�`������(p'N�yW�$��I��`����|�e@'��|�-r��䎴a�өÖ�G��r�[����͎&&֑�QD��|٠�2GRF|����σ���c�-\�-�E	xɽ��d~���u�&2�ن��͏�]k��ē��)ޤ8qE����!��0�]�K�~�?$M�R�;{[��b�O���RK�����׆*������T2�/��1�
�L8FR��J�sW_���^�gKYD��N��j̆D}XŌ���R�x]g��et���B��&]�uN�ڡ��t�β:9�?Jt#t�����e�����A4��_�B��F���n�7)G���]��L�{�Z�;��6��� KB--8}�D�+Μ� !ա9�����u����@�5�]��r��TZ��[L���ԫ㺯�7�IX"9I�Xyj�:~��fE�
�G�K���Q��H���ͩ7�m[}"�v��20w;M����;s%������i59�p� �����Pfw}�^{��7љ,���Xܗ��u��Y�/�=��xB�oLc��o�!Vc���G?�t>�;��K�V;���"^���P���̶Sjn�L����3�x�M�����][y%ٍyj�D��7lW��Z�9�V�ٱ��N�bl�j�牞yK��˄�^�rdv��AWzU�Ht1o�s��ʧ�n�Qi�)���<���B�!(5�a�W��2̓U�yw����D�a<�toa��s��4mF���Q�}f�MS0g��d�7�\�`ግ|i��ŋ��l���)M�|����h)�R<Y�SdDA��ՆK08�����h��|�EI������۩"�s&ʑ���U�M�-O��mNqb۾��JT�8�(ha���z�ِ����CG²��)(G��I ��������i�3д�9�����!��wD��f��׉`Db��6��<�n��t�B������D��ʈO_���*�lp����+���_�%����������\ل�3�3�	$���7I�P�wB�t/�j�om�������z�h���_�eٓ�>�9�7����;��}$���in�>t��ӧ-o�N!��T���o	�d1�X���s�0��w��;Ľ�a����S�0�n_����� ��)Ey��l6Fm~�h�d�a�%
f��OEm�}��h�����Z�������S&k&>�e=TB��u� ��l��x�f=p5�r�*�(V��*z��^Gv^�W��4��^-�����b;]��5��g��a��������D�s~
��D�e=�>V��w���࿎�K��W(���gWC�>Ƥ2�ݶ���$<B�T.�ҋgs剝�,Bd�{� ���1#���1�+�u����3fQWdIS�5��Q2XlD~�D�D$0$�L)-���Ji&��`Ir�$P�M%u˞
40�Z�%,��PL��9d5��4PW��<��*Ι��1�f�Pj�d�
���	��ҪR�⽘TY�5��Ff|x(+������Qv��2)`P�ȹ��Yi��Y�z��gK��l�����IV ���`���6̫0�V�e��_)�¨?����s��PzX�#�&)�:)sH$�˵(l�?>z�84�����cA�8��1���n������2@��ul�A����{��/�<TQB�'��>.��s�ze�v���*ny7